// DE0Qsys.v

// Generated using ACDS version 13.0sp1 232 at 2023.05.17.17:27:06

`timescale 1 ps / 1 ps
module DE0Qsys (
		input  wire        clk_50m_clk,           //        clk_50m.clk
		input  wire        reset_reset_n,         //          reset.reset_n
		output wire        dram_clk_clk,          //       dram_clk.clk
		input  wire        areset_export,         //         areset.export
		output wire        locked_export,         //         locked.export
		output wire        phasedone_export,      //      phasedone.export
		output wire [11:0] sdram_wires_addr,      //    sdram_wires.addr
		output wire [1:0]  sdram_wires_ba,        //               .ba
		output wire        sdram_wires_cas_n,     //               .cas_n
		output wire        sdram_wires_cke,       //               .cke
		output wire        sdram_wires_cs_n,      //               .cs_n
		inout  wire [15:0] sdram_wires_dq,        //               .dq
		output wire [1:0]  sdram_wires_dqm,       //               .dqm
		output wire        sdram_wires_ras_n,     //               .ras_n
		output wire        sdram_wires_we_n,      //               .we_n
		output wire [9:0]  led_export,            //            led.export
		input  wire [1:0]  button_export,         //         button.export
		input  wire [9:0]  sw_export,             //             sw.export
		output wire [7:0]  hex_0_export,          //          hex_0.export
		output wire [7:0]  motora_duty_export,    //    motora_duty.export
		output wire [7:0]  motorb_duty_export,    //    motorb_duty.export
		output wire [1:0]  motora_dir_export,     //     motora_dir.export
		output wire [1:0]  motorb_dir_export,     //     motorb_dir.export
		output wire [7:0]  hex_1_export,          //          hex_1.export
		input  wire        infra_sensor_0_export, // infra_sensor_0.export
		input  wire        infra_sensor_4_export, // infra_sensor_4.export
		input  wire        infra_sensor_3_export, // infra_sensor_3.export
		input  wire        infra_sensor_2_export, // infra_sensor_2.export
		input  wire        infra_sensor_1_export  // infra_sensor_1.export
	);

	wire          syspll_c0_clk;                                                                                    // syspll:c0 -> [APB:clk, APB_m0_translator:clk, APB_m0_translator_avalon_universal_master_0_agent:clk, APB_s0_translator:clk, APB_s0_translator_avalon_universal_slave_0_agent:clk, APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, crosser:in_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:in_clk, crosser_005:in_clk, crosser_006:in_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, crosser_010:in_clk, crosser_011:in_clk, crosser_012:in_clk, crosser_013:in_clk, crosser_014:in_clk, crosser_015:in_clk, crosser_016:in_clk, crosser_017:in_clk, crosser_018:out_clk, crosser_019:out_clk, crosser_020:out_clk, crosser_021:out_clk, crosser_022:out_clk, crosser_023:out_clk, crosser_024:out_clk, crosser_025:out_clk, crosser_026:out_clk, crosser_027:out_clk, crosser_028:out_clk, crosser_029:out_clk, crosser_030:out_clk, crosser_031:out_clk, crosser_032:out_clk, crosser_033:out_clk, dma:clk, dma_control_port_slave_translator:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_read_master_translator:clk, dma_read_master_translator_avalon_universal_master_0_agent:clk, dma_write_master_translator:clk, dma_write_master_translator_avalon_universal_master_0_agent:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_004:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, limiter:clk, limiter_001:clk, nios2cpu:clk, nios2cpu_data_master_translator:clk, nios2cpu_data_master_translator_avalon_universal_master_0_agent:clk, nios2cpu_instruction_master_translator:clk, nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2cpu_jtag_debug_module_translator:clk, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_004:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rsp_xbar_mux_003:clk, rsp_xbar_mux_004:clk, rst_controller:clk, sdram_ctrl:clk, sdram_ctrl_s1_translator:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	wire          syspll_c2_clk;                                                                                    // syspll:c2 -> [button:clk, button_s1_translator:clk, button_s1_translator_avalon_universal_slave_0_agent:clk, button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, crosser_002:out_clk, crosser_003:out_clk, crosser_004:out_clk, crosser_005:out_clk, crosser_006:out_clk, crosser_007:out_clk, crosser_008:out_clk, crosser_009:out_clk, crosser_010:out_clk, crosser_011:out_clk, crosser_012:out_clk, crosser_013:out_clk, crosser_014:out_clk, crosser_015:out_clk, crosser_016:out_clk, crosser_017:out_clk, crosser_018:in_clk, crosser_019:in_clk, crosser_020:in_clk, crosser_021:in_clk, crosser_022:in_clk, crosser_023:in_clk, crosser_024:in_clk, crosser_025:in_clk, crosser_026:in_clk, crosser_027:in_clk, crosser_028:in_clk, crosser_029:in_clk, crosser_030:in_clk, crosser_031:in_clk, crosser_032:in_clk, crosser_033:in_clk, hex_0:clk, hex_0_s1_translator:clk, hex_0_s1_translator_avalon_universal_slave_0_agent:clk, hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, hex_1:clk, hex_1_s1_translator:clk, hex_1_s1_translator_avalon_universal_slave_0_agent:clk, hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, infra_sensor_0:clk, infra_sensor_0_s1_translator:clk, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:clk, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, infra_sensor_1:clk, infra_sensor_1_s1_translator:clk, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:clk, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, infra_sensor_2:clk, infra_sensor_2_s1_translator:clk, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:clk, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, infra_sensor_3:clk, infra_sensor_3_s1_translator:clk, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:clk, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, infra_sensor_4:clk, infra_sensor_4_s1_translator:clk, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:clk, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led:clk, led_s1_translator:clk, led_s1_translator_avalon_universal_slave_0_agent:clk, led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, motorA_dir:clk, motorA_dir_s1_translator:clk, motorA_dir_s1_translator_avalon_universal_slave_0_agent:clk, motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, motorA_duty:clk, motorA_duty_s1_translator:clk, motorA_duty_s1_translator_avalon_universal_slave_0_agent:clk, motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, motorB_dir:clk, motorB_dir_s1_translator:clk, motorB_dir_s1_translator_avalon_universal_slave_0_agent:clk, motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, motorB_duty:clk, motorB_duty_s1_translator:clk, motorB_duty_s1_translator_avalon_universal_slave_0_agent:clk, motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rst_controller_001:clk, sw:clk, sw_s1_translator:clk, sw_s1_translator_avalon_universal_slave_0_agent:clk, sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire          nios2cpu_instruction_master_waitrequest;                                                          // nios2cpu_instruction_master_translator:av_waitrequest -> nios2cpu:i_waitrequest
	wire   [25:0] nios2cpu_instruction_master_address;                                                              // nios2cpu:i_address -> nios2cpu_instruction_master_translator:av_address
	wire          nios2cpu_instruction_master_read;                                                                 // nios2cpu:i_read -> nios2cpu_instruction_master_translator:av_read
	wire   [31:0] nios2cpu_instruction_master_readdata;                                                             // nios2cpu_instruction_master_translator:av_readdata -> nios2cpu:i_readdata
	wire          nios2cpu_data_master_waitrequest;                                                                 // nios2cpu_data_master_translator:av_waitrequest -> nios2cpu:d_waitrequest
	wire   [31:0] nios2cpu_data_master_writedata;                                                                   // nios2cpu:d_writedata -> nios2cpu_data_master_translator:av_writedata
	wire   [25:0] nios2cpu_data_master_address;                                                                     // nios2cpu:d_address -> nios2cpu_data_master_translator:av_address
	wire          nios2cpu_data_master_write;                                                                       // nios2cpu:d_write -> nios2cpu_data_master_translator:av_write
	wire          nios2cpu_data_master_read;                                                                        // nios2cpu:d_read -> nios2cpu_data_master_translator:av_read
	wire   [31:0] nios2cpu_data_master_readdata;                                                                    // nios2cpu_data_master_translator:av_readdata -> nios2cpu:d_readdata
	wire          nios2cpu_data_master_debugaccess;                                                                 // nios2cpu:jtag_debug_module_debugaccess_to_roms -> nios2cpu_data_master_translator:av_debugaccess
	wire    [3:0] nios2cpu_data_master_byteenable;                                                                  // nios2cpu:d_byteenable -> nios2cpu_data_master_translator:av_byteenable
	wire    [7:0] dma_read_master_burstcount;                                                                       // dma:read_burstcount -> dma_read_master_translator:av_burstcount
	wire          dma_read_master_waitrequest;                                                                      // dma_read_master_translator:av_waitrequest -> dma:read_waitrequest
	wire   [25:0] dma_read_master_address;                                                                          // dma:read_address -> dma_read_master_translator:av_address
	wire          dma_read_master_chipselect;                                                                       // dma:read_chipselect -> dma_read_master_translator:av_chipselect
	wire          dma_read_master_read;                                                                             // dma:read_read_n -> dma_read_master_translator:av_read
	wire   [31:0] dma_read_master_readdata;                                                                         // dma_read_master_translator:av_readdata -> dma:read_readdata
	wire          dma_read_master_readdatavalid;                                                                    // dma_read_master_translator:av_readdatavalid -> dma:read_readdatavalid
	wire    [7:0] dma_write_master_burstcount;                                                                      // dma:write_burstcount -> dma_write_master_translator:av_burstcount
	wire          dma_write_master_waitrequest;                                                                     // dma_write_master_translator:av_waitrequest -> dma:write_waitrequest
	wire   [31:0] dma_write_master_writedata;                                                                       // dma:write_writedata -> dma_write_master_translator:av_writedata
	wire   [25:0] dma_write_master_address;                                                                         // dma:write_address -> dma_write_master_translator:av_address
	wire          dma_write_master_chipselect;                                                                      // dma:write_chipselect -> dma_write_master_translator:av_chipselect
	wire          dma_write_master_write;                                                                           // dma:write_write_n -> dma_write_master_translator:av_write
	wire    [3:0] dma_write_master_byteenable;                                                                      // dma:write_byteenable -> dma_write_master_translator:av_byteenable
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                            // nios2cpu:jtag_debug_module_waitrequest -> nios2cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                              // nios2cpu_jtag_debug_module_translator:av_writedata -> nios2cpu:jtag_debug_module_writedata
	wire    [8:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                // nios2cpu_jtag_debug_module_translator:av_address -> nios2cpu:jtag_debug_module_address
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                  // nios2cpu_jtag_debug_module_translator:av_write -> nios2cpu:jtag_debug_module_write
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                   // nios2cpu_jtag_debug_module_translator:av_read -> nios2cpu:jtag_debug_module_read
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                               // nios2cpu:jtag_debug_module_readdata -> nios2cpu_jtag_debug_module_translator:av_readdata
	wire          nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                            // nios2cpu_jtag_debug_module_translator:av_debugaccess -> nios2cpu:jtag_debug_module_debugaccess
	wire    [3:0] nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                             // nios2cpu_jtag_debug_module_translator:av_byteenable -> nios2cpu:jtag_debug_module_byteenable
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest;                                         // sdram_ctrl:za_waitrequest -> sdram_ctrl_s1_translator:av_waitrequest
	wire   [15:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata;                                           // sdram_ctrl_s1_translator:av_writedata -> sdram_ctrl:az_data
	wire   [21:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_address;                                             // sdram_ctrl_s1_translator:av_address -> sdram_ctrl:az_addr
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect;                                          // sdram_ctrl_s1_translator:av_chipselect -> sdram_ctrl:az_cs
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_write;                                               // sdram_ctrl_s1_translator:av_write -> sdram_ctrl:az_wr_n
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_read;                                                // sdram_ctrl_s1_translator:av_read -> sdram_ctrl:az_rd_n
	wire   [15:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata;                                            // sdram_ctrl:za_data -> sdram_ctrl_s1_translator:av_readdata
	wire          sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid;                                       // sdram_ctrl:za_valid -> sdram_ctrl_s1_translator:av_readdatavalid
	wire    [1:0] sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable;                                          // sdram_ctrl_s1_translator:av_byteenable -> sdram_ctrl:az_be_n
	wire          apb_s0_translator_avalon_anti_slave_0_waitrequest;                                                // APB:s0_waitrequest -> APB_s0_translator:av_waitrequest
	wire    [0:0] apb_s0_translator_avalon_anti_slave_0_burstcount;                                                 // APB_s0_translator:av_burstcount -> APB:s0_burstcount
	wire   [31:0] apb_s0_translator_avalon_anti_slave_0_writedata;                                                  // APB_s0_translator:av_writedata -> APB:s0_writedata
	wire    [9:0] apb_s0_translator_avalon_anti_slave_0_address;                                                    // APB_s0_translator:av_address -> APB:s0_address
	wire          apb_s0_translator_avalon_anti_slave_0_write;                                                      // APB_s0_translator:av_write -> APB:s0_write
	wire          apb_s0_translator_avalon_anti_slave_0_read;                                                       // APB_s0_translator:av_read -> APB:s0_read
	wire   [31:0] apb_s0_translator_avalon_anti_slave_0_readdata;                                                   // APB:s0_readdata -> APB_s0_translator:av_readdata
	wire          apb_s0_translator_avalon_anti_slave_0_debugaccess;                                                // APB_s0_translator:av_debugaccess -> APB:s0_debugaccess
	wire          apb_s0_translator_avalon_anti_slave_0_readdatavalid;                                              // APB:s0_readdatavalid -> APB_s0_translator:av_readdatavalid
	wire    [3:0] apb_s0_translator_avalon_anti_slave_0_byteenable;                                                 // APB_s0_translator:av_byteenable -> APB:s0_byteenable
	wire   [31:0] syspll_pll_slave_translator_avalon_anti_slave_0_writedata;                                        // syspll_pll_slave_translator:av_writedata -> syspll:writedata
	wire    [1:0] syspll_pll_slave_translator_avalon_anti_slave_0_address;                                          // syspll_pll_slave_translator:av_address -> syspll:address
	wire          syspll_pll_slave_translator_avalon_anti_slave_0_write;                                            // syspll_pll_slave_translator:av_write -> syspll:write
	wire          syspll_pll_slave_translator_avalon_anti_slave_0_read;                                             // syspll_pll_slave_translator:av_read -> syspll:read
	wire   [31:0] syspll_pll_slave_translator_avalon_anti_slave_0_readdata;                                         // syspll:readdata -> syspll_pll_slave_translator:av_readdata
	wire   [25:0] dma_control_port_slave_translator_avalon_anti_slave_0_writedata;                                  // dma_control_port_slave_translator:av_writedata -> dma:dma_ctl_writedata
	wire    [2:0] dma_control_port_slave_translator_avalon_anti_slave_0_address;                                    // dma_control_port_slave_translator:av_address -> dma:dma_ctl_address
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                 // dma_control_port_slave_translator:av_chipselect -> dma:dma_ctl_chipselect
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_write;                                      // dma_control_port_slave_translator:av_write -> dma:dma_ctl_write_n
	wire   [25:0] dma_control_port_slave_translator_avalon_anti_slave_0_readdata;                                   // dma:dma_ctl_readdata -> dma_control_port_slave_translator:av_readdata
	wire    [0:0] apb_m0_burstcount;                                                                                // APB:m0_burstcount -> APB_m0_translator:av_burstcount
	wire          apb_m0_waitrequest;                                                                               // APB_m0_translator:av_waitrequest -> APB:m0_waitrequest
	wire    [9:0] apb_m0_address;                                                                                   // APB:m0_address -> APB_m0_translator:av_address
	wire   [31:0] apb_m0_writedata;                                                                                 // APB:m0_writedata -> APB_m0_translator:av_writedata
	wire          apb_m0_write;                                                                                     // APB:m0_write -> APB_m0_translator:av_write
	wire          apb_m0_read;                                                                                      // APB:m0_read -> APB_m0_translator:av_read
	wire   [31:0] apb_m0_readdata;                                                                                  // APB_m0_translator:av_readdata -> APB:m0_readdata
	wire          apb_m0_debugaccess;                                                                               // APB:m0_debugaccess -> APB_m0_translator:av_debugaccess
	wire    [3:0] apb_m0_byteenable;                                                                                // APB:m0_byteenable -> APB_m0_translator:av_byteenable
	wire          apb_m0_readdatavalid;                                                                             // APB_m0_translator:av_readdatavalid -> APB:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                  // led_s1_translator:av_writedata -> led:writedata
	wire    [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                    // led_s1_translator:av_address -> led:address
	wire          led_s1_translator_avalon_anti_slave_0_chipselect;                                                 // led_s1_translator:av_chipselect -> led:chipselect
	wire          led_s1_translator_avalon_anti_slave_0_write;                                                      // led_s1_translator:av_write -> led:write_n
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                   // led:readdata -> led_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                  // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                    // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer:readdata -> timer_s1_translator:av_readdata
	wire   [31:0] button_s1_translator_avalon_anti_slave_0_writedata;                                               // button_s1_translator:av_writedata -> button:writedata
	wire    [1:0] button_s1_translator_avalon_anti_slave_0_address;                                                 // button_s1_translator:av_address -> button:address
	wire          button_s1_translator_avalon_anti_slave_0_chipselect;                                              // button_s1_translator:av_chipselect -> button:chipselect
	wire          button_s1_translator_avalon_anti_slave_0_write;                                                   // button_s1_translator:av_write -> button:write_n
	wire   [31:0] button_s1_translator_avalon_anti_slave_0_readdata;                                                // button:readdata -> button_s1_translator:av_readdata
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_writedata;                                                   // sw_s1_translator:av_writedata -> sw:writedata
	wire    [1:0] sw_s1_translator_avalon_anti_slave_0_address;                                                     // sw_s1_translator:av_address -> sw:address
	wire          sw_s1_translator_avalon_anti_slave_0_chipselect;                                                  // sw_s1_translator:av_chipselect -> sw:chipselect
	wire          sw_s1_translator_avalon_anti_slave_0_write;                                                       // sw_s1_translator:av_write -> sw:write_n
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_readdata;                                                    // sw:readdata -> sw_s1_translator:av_readdata
	wire   [31:0] hex_0_s1_translator_avalon_anti_slave_0_writedata;                                                // hex_0_s1_translator:av_writedata -> hex_0:writedata
	wire    [1:0] hex_0_s1_translator_avalon_anti_slave_0_address;                                                  // hex_0_s1_translator:av_address -> hex_0:address
	wire          hex_0_s1_translator_avalon_anti_slave_0_chipselect;                                               // hex_0_s1_translator:av_chipselect -> hex_0:chipselect
	wire          hex_0_s1_translator_avalon_anti_slave_0_write;                                                    // hex_0_s1_translator:av_write -> hex_0:write_n
	wire   [31:0] hex_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // hex_0:readdata -> hex_0_s1_translator:av_readdata
	wire   [31:0] motora_duty_s1_translator_avalon_anti_slave_0_writedata;                                          // motorA_duty_s1_translator:av_writedata -> motorA_duty:writedata
	wire    [1:0] motora_duty_s1_translator_avalon_anti_slave_0_address;                                            // motorA_duty_s1_translator:av_address -> motorA_duty:address
	wire          motora_duty_s1_translator_avalon_anti_slave_0_chipselect;                                         // motorA_duty_s1_translator:av_chipselect -> motorA_duty:chipselect
	wire          motora_duty_s1_translator_avalon_anti_slave_0_write;                                              // motorA_duty_s1_translator:av_write -> motorA_duty:write_n
	wire   [31:0] motora_duty_s1_translator_avalon_anti_slave_0_readdata;                                           // motorA_duty:readdata -> motorA_duty_s1_translator:av_readdata
	wire   [31:0] motorb_duty_s1_translator_avalon_anti_slave_0_writedata;                                          // motorB_duty_s1_translator:av_writedata -> motorB_duty:writedata
	wire    [1:0] motorb_duty_s1_translator_avalon_anti_slave_0_address;                                            // motorB_duty_s1_translator:av_address -> motorB_duty:address
	wire          motorb_duty_s1_translator_avalon_anti_slave_0_chipselect;                                         // motorB_duty_s1_translator:av_chipselect -> motorB_duty:chipselect
	wire          motorb_duty_s1_translator_avalon_anti_slave_0_write;                                              // motorB_duty_s1_translator:av_write -> motorB_duty:write_n
	wire   [31:0] motorb_duty_s1_translator_avalon_anti_slave_0_readdata;                                           // motorB_duty:readdata -> motorB_duty_s1_translator:av_readdata
	wire   [31:0] motora_dir_s1_translator_avalon_anti_slave_0_writedata;                                           // motorA_dir_s1_translator:av_writedata -> motorA_dir:writedata
	wire    [1:0] motora_dir_s1_translator_avalon_anti_slave_0_address;                                             // motorA_dir_s1_translator:av_address -> motorA_dir:address
	wire          motora_dir_s1_translator_avalon_anti_slave_0_chipselect;                                          // motorA_dir_s1_translator:av_chipselect -> motorA_dir:chipselect
	wire          motora_dir_s1_translator_avalon_anti_slave_0_write;                                               // motorA_dir_s1_translator:av_write -> motorA_dir:write_n
	wire   [31:0] motora_dir_s1_translator_avalon_anti_slave_0_readdata;                                            // motorA_dir:readdata -> motorA_dir_s1_translator:av_readdata
	wire   [31:0] motorb_dir_s1_translator_avalon_anti_slave_0_writedata;                                           // motorB_dir_s1_translator:av_writedata -> motorB_dir:writedata
	wire    [1:0] motorb_dir_s1_translator_avalon_anti_slave_0_address;                                             // motorB_dir_s1_translator:av_address -> motorB_dir:address
	wire          motorb_dir_s1_translator_avalon_anti_slave_0_chipselect;                                          // motorB_dir_s1_translator:av_chipselect -> motorB_dir:chipselect
	wire          motorb_dir_s1_translator_avalon_anti_slave_0_write;                                               // motorB_dir_s1_translator:av_write -> motorB_dir:write_n
	wire   [31:0] motorb_dir_s1_translator_avalon_anti_slave_0_readdata;                                            // motorB_dir:readdata -> motorB_dir_s1_translator:av_readdata
	wire   [31:0] hex_1_s1_translator_avalon_anti_slave_0_writedata;                                                // hex_1_s1_translator:av_writedata -> hex_1:writedata
	wire    [1:0] hex_1_s1_translator_avalon_anti_slave_0_address;                                                  // hex_1_s1_translator:av_address -> hex_1:address
	wire          hex_1_s1_translator_avalon_anti_slave_0_chipselect;                                               // hex_1_s1_translator:av_chipselect -> hex_1:chipselect
	wire          hex_1_s1_translator_avalon_anti_slave_0_write;                                                    // hex_1_s1_translator:av_write -> hex_1:write_n
	wire   [31:0] hex_1_s1_translator_avalon_anti_slave_0_readdata;                                                 // hex_1:readdata -> hex_1_s1_translator:av_readdata
	wire    [1:0] infra_sensor_0_s1_translator_avalon_anti_slave_0_address;                                         // infra_sensor_0_s1_translator:av_address -> infra_sensor_0:address
	wire   [31:0] infra_sensor_0_s1_translator_avalon_anti_slave_0_readdata;                                        // infra_sensor_0:readdata -> infra_sensor_0_s1_translator:av_readdata
	wire    [1:0] infra_sensor_1_s1_translator_avalon_anti_slave_0_address;                                         // infra_sensor_1_s1_translator:av_address -> infra_sensor_1:address
	wire   [31:0] infra_sensor_1_s1_translator_avalon_anti_slave_0_readdata;                                        // infra_sensor_1:readdata -> infra_sensor_1_s1_translator:av_readdata
	wire    [1:0] infra_sensor_2_s1_translator_avalon_anti_slave_0_address;                                         // infra_sensor_2_s1_translator:av_address -> infra_sensor_2:address
	wire   [31:0] infra_sensor_2_s1_translator_avalon_anti_slave_0_readdata;                                        // infra_sensor_2:readdata -> infra_sensor_2_s1_translator:av_readdata
	wire    [1:0] infra_sensor_3_s1_translator_avalon_anti_slave_0_address;                                         // infra_sensor_3_s1_translator:av_address -> infra_sensor_3:address
	wire   [31:0] infra_sensor_3_s1_translator_avalon_anti_slave_0_readdata;                                        // infra_sensor_3:readdata -> infra_sensor_3_s1_translator:av_readdata
	wire    [1:0] infra_sensor_4_s1_translator_avalon_anti_slave_0_address;                                         // infra_sensor_4_s1_translator:av_address -> infra_sensor_4:address
	wire   [31:0] infra_sensor_4_s1_translator_avalon_anti_slave_0_readdata;                                        // infra_sensor_4:readdata -> infra_sensor_4_s1_translator:av_readdata
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                     // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                      // nios2cpu_instruction_master_translator:uav_burstcount -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata;                       // nios2cpu_instruction_master_translator:uav_writedata -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_address;                         // nios2cpu_instruction_master_translator:uav_address -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_lock;                            // nios2cpu_instruction_master_translator:uav_lock -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_write;                           // nios2cpu_instruction_master_translator:uav_write -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_read;                            // nios2cpu_instruction_master_translator:uav_read -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata;                        // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2cpu_instruction_master_translator:uav_readdata
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                     // nios2cpu_instruction_master_translator:uav_debugaccess -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                      // nios2cpu_instruction_master_translator:uav_byteenable -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                   // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2cpu_instruction_master_translator:uav_readdatavalid
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest;                            // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2cpu_data_master_translator:uav_waitrequest
	wire    [2:0] nios2cpu_data_master_translator_avalon_universal_master_0_burstcount;                             // nios2cpu_data_master_translator:uav_burstcount -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2cpu_data_master_translator_avalon_universal_master_0_writedata;                              // nios2cpu_data_master_translator:uav_writedata -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2cpu_data_master_translator_avalon_universal_master_0_address;                                // nios2cpu_data_master_translator:uav_address -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_lock;                                   // nios2cpu_data_master_translator:uav_lock -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_write;                                  // nios2cpu_data_master_translator:uav_write -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_read;                                   // nios2cpu_data_master_translator:uav_read -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2cpu_data_master_translator_avalon_universal_master_0_readdata;                               // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2cpu_data_master_translator:uav_readdata
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess;                            // nios2cpu_data_master_translator:uav_debugaccess -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2cpu_data_master_translator_avalon_universal_master_0_byteenable;                             // nios2cpu_data_master_translator:uav_byteenable -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                          // nios2cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2cpu_data_master_translator:uav_readdatavalid
	wire          dma_read_master_translator_avalon_universal_master_0_waitrequest;                                 // dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_read_master_translator:uav_waitrequest
	wire    [9:0] dma_read_master_translator_avalon_universal_master_0_burstcount;                                  // dma_read_master_translator:uav_burstcount -> dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_writedata;                                   // dma_read_master_translator:uav_writedata -> dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] dma_read_master_translator_avalon_universal_master_0_address;                                     // dma_read_master_translator:uav_address -> dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_read_master_translator_avalon_universal_master_0_lock;                                        // dma_read_master_translator:uav_lock -> dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_read_master_translator_avalon_universal_master_0_write;                                       // dma_read_master_translator:uav_write -> dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_read_master_translator_avalon_universal_master_0_read;                                        // dma_read_master_translator:uav_read -> dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_readdata;                                    // dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_read_master_translator:uav_readdata
	wire          dma_read_master_translator_avalon_universal_master_0_debugaccess;                                 // dma_read_master_translator:uav_debugaccess -> dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_read_master_translator_avalon_universal_master_0_byteenable;                                  // dma_read_master_translator:uav_byteenable -> dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_read_master_translator_avalon_universal_master_0_readdatavalid;                               // dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_read_master_translator:uav_readdatavalid
	wire          dma_write_master_translator_avalon_universal_master_0_waitrequest;                                // dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_write_master_translator:uav_waitrequest
	wire    [9:0] dma_write_master_translator_avalon_universal_master_0_burstcount;                                 // dma_write_master_translator:uav_burstcount -> dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_writedata;                                  // dma_write_master_translator:uav_writedata -> dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] dma_write_master_translator_avalon_universal_master_0_address;                                    // dma_write_master_translator:uav_address -> dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_write_master_translator_avalon_universal_master_0_lock;                                       // dma_write_master_translator:uav_lock -> dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_write_master_translator_avalon_universal_master_0_write;                                      // dma_write_master_translator:uav_write -> dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_write_master_translator_avalon_universal_master_0_read;                                       // dma_write_master_translator:uav_read -> dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_readdata;                                   // dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_write_master_translator:uav_readdata
	wire          dma_write_master_translator_avalon_universal_master_0_debugaccess;                                // dma_write_master_translator:uav_debugaccess -> dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_write_master_translator_avalon_universal_master_0_byteenable;                                 // dma_write_master_translator:uav_byteenable -> dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_write_master_translator_avalon_universal_master_0_readdatavalid;                              // dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_write_master_translator:uav_readdatavalid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // nios2cpu_jtag_debug_module_translator:uav_waitrequest -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;               // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2cpu_jtag_debug_module_translator:uav_writedata
	wire   [25:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                  // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2cpu_jtag_debug_module_translator:uav_address
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2cpu_jtag_debug_module_translator:uav_write
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2cpu_jtag_debug_module_translator:uav_lock
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                 // nios2cpu_jtag_debug_module_translator:uav_readdata -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // nios2cpu_jtag_debug_module_translator:uav_readdatavalid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;               // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2cpu_jtag_debug_module_translator:uav_byteenable
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;             // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;             // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // sdram_ctrl_s1_translator:uav_waitrequest -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_ctrl_s1_translator:uav_burstcount
	wire   [15:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_ctrl_s1_translator:uav_writedata
	wire   [25:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_ctrl_s1_translator:uav_address
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_ctrl_s1_translator:uav_write
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_ctrl_s1_translator:uav_lock
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_ctrl_s1_translator:uav_read
	wire   [15:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // sdram_ctrl_s1_translator:uav_readdata -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // sdram_ctrl_s1_translator:uav_readdatavalid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_ctrl_s1_translator:uav_debugaccess
	wire    [1:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_ctrl_s1_translator:uav_byteenable
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [88:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [88:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // APB_s0_translator:uav_waitrequest -> APB_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // APB_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> APB_s0_translator:uav_burstcount
	wire   [31:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // APB_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> APB_s0_translator:uav_writedata
	wire   [25:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_address;                                      // APB_s0_translator_avalon_universal_slave_0_agent:m0_address -> APB_s0_translator:uav_address
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_write;                                        // APB_s0_translator_avalon_universal_slave_0_agent:m0_write -> APB_s0_translator:uav_write
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                         // APB_s0_translator_avalon_universal_slave_0_agent:m0_lock -> APB_s0_translator:uav_lock
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_read;                                         // APB_s0_translator_avalon_universal_slave_0_agent:m0_read -> APB_s0_translator:uav_read
	wire   [31:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // APB_s0_translator:uav_readdata -> APB_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // APB_s0_translator:uav_readdatavalid -> APB_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // APB_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> APB_s0_translator:uav_debugaccess
	wire    [3:0] apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // APB_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> APB_s0_translator:uav_byteenable
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // APB_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // APB_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // syspll_pll_slave_translator:uav_waitrequest -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> syspll_pll_slave_translator:uav_burstcount
	wire   [31:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> syspll_pll_slave_translator:uav_writedata
	wire   [25:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> syspll_pll_slave_translator:uav_address
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> syspll_pll_slave_translator:uav_write
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> syspll_pll_slave_translator:uav_lock
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> syspll_pll_slave_translator:uav_read
	wire   [31:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // syspll_pll_slave_translator:uav_readdata -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // syspll_pll_slave_translator:uav_readdatavalid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> syspll_pll_slave_translator:uav_debugaccess
	wire    [3:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // syspll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> syspll_pll_slave_translator:uav_byteenable
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // dma_control_port_slave_translator:uav_waitrequest -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_control_port_slave_translator:uav_writedata
	wire   [25:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_control_port_slave_translator:uav_address
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_control_port_slave_translator:uav_write
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_control_port_slave_translator:uav_lock
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_control_port_slave_translator:uav_read
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // dma_control_port_slave_translator:uav_readdata -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // dma_control_port_slave_translator:uav_readdatavalid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_control_port_slave_translator:uav_byteenable
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          apb_m0_translator_avalon_universal_master_0_waitrequest;                                          // APB_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> APB_m0_translator:uav_waitrequest
	wire    [2:0] apb_m0_translator_avalon_universal_master_0_burstcount;                                           // APB_m0_translator:uav_burstcount -> APB_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] apb_m0_translator_avalon_universal_master_0_writedata;                                            // APB_m0_translator:uav_writedata -> APB_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] apb_m0_translator_avalon_universal_master_0_address;                                              // APB_m0_translator:uav_address -> APB_m0_translator_avalon_universal_master_0_agent:av_address
	wire          apb_m0_translator_avalon_universal_master_0_lock;                                                 // APB_m0_translator:uav_lock -> APB_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          apb_m0_translator_avalon_universal_master_0_write;                                                // APB_m0_translator:uav_write -> APB_m0_translator_avalon_universal_master_0_agent:av_write
	wire          apb_m0_translator_avalon_universal_master_0_read;                                                 // APB_m0_translator:uav_read -> APB_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] apb_m0_translator_avalon_universal_master_0_readdata;                                             // APB_m0_translator_avalon_universal_master_0_agent:av_readdata -> APB_m0_translator:uav_readdata
	wire          apb_m0_translator_avalon_universal_master_0_debugaccess;                                          // APB_m0_translator:uav_debugaccess -> APB_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] apb_m0_translator_avalon_universal_master_0_byteenable;                                           // APB_m0_translator:uav_byteenable -> APB_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          apb_m0_translator_avalon_universal_master_0_readdatavalid;                                        // APB_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> APB_m0_translator:uav_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire    [9:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire    [9:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire    [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire    [9:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // button_s1_translator:uav_waitrequest -> button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_s1_translator:uav_burstcount
	wire   [31:0] button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_s1_translator:uav_writedata
	wire    [9:0] button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // button_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_s1_translator:uav_address
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // button_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_s1_translator:uav_write
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_s1_translator:uav_lock
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // button_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_s1_translator:uav_read
	wire   [31:0] button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // button_s1_translator:uav_readdata -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // button_s1_translator:uav_readdatavalid -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_s1_translator:uav_debugaccess
	wire    [3:0] button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_s1_translator:uav_byteenable
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sw_s1_translator:uav_waitrequest -> sw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sw_s1_translator:uav_burstcount
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sw_s1_translator:uav_writedata
	wire    [9:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // sw_s1_translator_avalon_universal_slave_0_agent:m0_address -> sw_s1_translator:uav_address
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // sw_s1_translator_avalon_universal_slave_0_agent:m0_write -> sw_s1_translator:uav_write
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sw_s1_translator:uav_lock
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // sw_s1_translator_avalon_universal_slave_0_agent:m0_read -> sw_s1_translator:uav_read
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sw_s1_translator:uav_readdata -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sw_s1_translator:uav_readdatavalid -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sw_s1_translator:uav_debugaccess
	wire    [3:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sw_s1_translator:uav_byteenable
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                             // sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                              // sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                             // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // hex_0_s1_translator:uav_waitrequest -> hex_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex_0_s1_translator:uav_burstcount
	wire   [31:0] hex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex_0_s1_translator:uav_writedata
	wire    [9:0] hex_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex_0_s1_translator:uav_address
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex_0_s1_translator:uav_write
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex_0_s1_translator:uav_lock
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex_0_s1_translator:uav_read
	wire   [31:0] hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // hex_0_s1_translator:uav_readdata -> hex_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // hex_0_s1_translator:uav_readdatavalid -> hex_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex_0_s1_translator:uav_debugaccess
	wire    [3:0] hex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // hex_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex_0_s1_translator:uav_byteenable
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // hex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // hex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // hex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // hex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // hex_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // hex_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // motorA_duty_s1_translator:uav_waitrequest -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motorA_duty_s1_translator:uav_burstcount
	wire   [31:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motorA_duty_s1_translator:uav_writedata
	wire    [9:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_address -> motorA_duty_s1_translator:uav_address
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_write -> motorA_duty_s1_translator:uav_write
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motorA_duty_s1_translator:uav_lock
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_read -> motorA_duty_s1_translator:uav_read
	wire   [31:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // motorA_duty_s1_translator:uav_readdata -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // motorA_duty_s1_translator:uav_readdatavalid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motorA_duty_s1_translator:uav_debugaccess
	wire    [3:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // motorA_duty_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motorA_duty_s1_translator:uav_byteenable
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // motorB_duty_s1_translator:uav_waitrequest -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motorB_duty_s1_translator:uav_burstcount
	wire   [31:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motorB_duty_s1_translator:uav_writedata
	wire    [9:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_address -> motorB_duty_s1_translator:uav_address
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_write -> motorB_duty_s1_translator:uav_write
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motorB_duty_s1_translator:uav_lock
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_read -> motorB_duty_s1_translator:uav_read
	wire   [31:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // motorB_duty_s1_translator:uav_readdata -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // motorB_duty_s1_translator:uav_readdatavalid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motorB_duty_s1_translator:uav_debugaccess
	wire    [3:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // motorB_duty_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motorB_duty_s1_translator:uav_byteenable
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // motorA_dir_s1_translator:uav_waitrequest -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motorA_dir_s1_translator:uav_burstcount
	wire   [31:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motorA_dir_s1_translator:uav_writedata
	wire    [9:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_address -> motorA_dir_s1_translator:uav_address
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_write -> motorA_dir_s1_translator:uav_write
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motorA_dir_s1_translator:uav_lock
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_read -> motorA_dir_s1_translator:uav_read
	wire   [31:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // motorA_dir_s1_translator:uav_readdata -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // motorA_dir_s1_translator:uav_readdatavalid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motorA_dir_s1_translator:uav_debugaccess
	wire    [3:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // motorA_dir_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motorA_dir_s1_translator:uav_byteenable
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // motorB_dir_s1_translator:uav_waitrequest -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motorB_dir_s1_translator:uav_burstcount
	wire   [31:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motorB_dir_s1_translator:uav_writedata
	wire    [9:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_address -> motorB_dir_s1_translator:uav_address
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_write -> motorB_dir_s1_translator:uav_write
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motorB_dir_s1_translator:uav_lock
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_read -> motorB_dir_s1_translator:uav_read
	wire   [31:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // motorB_dir_s1_translator:uav_readdata -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // motorB_dir_s1_translator:uav_readdatavalid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motorB_dir_s1_translator:uav_debugaccess
	wire    [3:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // motorB_dir_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motorB_dir_s1_translator:uav_byteenable
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // hex_1_s1_translator:uav_waitrequest -> hex_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex_1_s1_translator:uav_burstcount
	wire   [31:0] hex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex_1_s1_translator:uav_writedata
	wire    [9:0] hex_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex_1_s1_translator:uav_address
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex_1_s1_translator:uav_write
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex_1_s1_translator:uav_lock
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex_1_s1_translator:uav_read
	wire   [31:0] hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // hex_1_s1_translator:uav_readdata -> hex_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // hex_1_s1_translator:uav_readdatavalid -> hex_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex_1_s1_translator:uav_debugaccess
	wire    [3:0] hex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // hex_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex_1_s1_translator:uav_byteenable
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // hex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // hex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // hex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // hex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // hex_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // hex_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // infra_sensor_0_s1_translator:uav_waitrequest -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> infra_sensor_0_s1_translator:uav_burstcount
	wire   [31:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> infra_sensor_0_s1_translator:uav_writedata
	wire    [9:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> infra_sensor_0_s1_translator:uav_address
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> infra_sensor_0_s1_translator:uav_write
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> infra_sensor_0_s1_translator:uav_lock
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> infra_sensor_0_s1_translator:uav_read
	wire   [31:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // infra_sensor_0_s1_translator:uav_readdata -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // infra_sensor_0_s1_translator:uav_readdatavalid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> infra_sensor_0_s1_translator:uav_debugaccess
	wire    [3:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> infra_sensor_0_s1_translator:uav_byteenable
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // infra_sensor_1_s1_translator:uav_waitrequest -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> infra_sensor_1_s1_translator:uav_burstcount
	wire   [31:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> infra_sensor_1_s1_translator:uav_writedata
	wire    [9:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> infra_sensor_1_s1_translator:uav_address
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> infra_sensor_1_s1_translator:uav_write
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> infra_sensor_1_s1_translator:uav_lock
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> infra_sensor_1_s1_translator:uav_read
	wire   [31:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // infra_sensor_1_s1_translator:uav_readdata -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // infra_sensor_1_s1_translator:uav_readdatavalid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> infra_sensor_1_s1_translator:uav_debugaccess
	wire    [3:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> infra_sensor_1_s1_translator:uav_byteenable
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // infra_sensor_2_s1_translator:uav_waitrequest -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> infra_sensor_2_s1_translator:uav_burstcount
	wire   [31:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> infra_sensor_2_s1_translator:uav_writedata
	wire    [9:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> infra_sensor_2_s1_translator:uav_address
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> infra_sensor_2_s1_translator:uav_write
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> infra_sensor_2_s1_translator:uav_lock
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> infra_sensor_2_s1_translator:uav_read
	wire   [31:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // infra_sensor_2_s1_translator:uav_readdata -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // infra_sensor_2_s1_translator:uav_readdatavalid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> infra_sensor_2_s1_translator:uav_debugaccess
	wire    [3:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> infra_sensor_2_s1_translator:uav_byteenable
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // infra_sensor_3_s1_translator:uav_waitrequest -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> infra_sensor_3_s1_translator:uav_burstcount
	wire   [31:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> infra_sensor_3_s1_translator:uav_writedata
	wire    [9:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> infra_sensor_3_s1_translator:uav_address
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> infra_sensor_3_s1_translator:uav_write
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> infra_sensor_3_s1_translator:uav_lock
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> infra_sensor_3_s1_translator:uav_read
	wire   [31:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // infra_sensor_3_s1_translator:uav_readdata -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // infra_sensor_3_s1_translator:uav_readdatavalid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> infra_sensor_3_s1_translator:uav_debugaccess
	wire    [3:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> infra_sensor_3_s1_translator:uav_byteenable
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // infra_sensor_4_s1_translator:uav_waitrequest -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> infra_sensor_4_s1_translator:uav_burstcount
	wire   [31:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> infra_sensor_4_s1_translator:uav_writedata
	wire    [9:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> infra_sensor_4_s1_translator:uav_address
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> infra_sensor_4_s1_translator:uav_write
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> infra_sensor_4_s1_translator:uav_lock
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> infra_sensor_4_s1_translator:uav_read
	wire   [31:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // infra_sensor_4_s1_translator:uav_readdata -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // infra_sensor_4_s1_translator:uav_readdatavalid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> infra_sensor_4_s1_translator:uav_debugaccess
	wire    [3:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> infra_sensor_4_s1_translator:uav_byteenable
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;            // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                  // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;          // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [105:0] nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                   // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router:sink_ready -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                         // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [105:0] nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                          // nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_001:sink_ready -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                              // dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [105:0] dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                               // dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_002:sink_ready -> dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                             // dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [105:0] dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                              // dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_003:sink_ready -> dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                    // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [105:0] nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                     // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [87:0] sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // APB_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                        // APB_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // APB_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [105:0] apb_s0_translator_avalon_universal_slave_0_agent_rp_data;                                         // APB_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          apb_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_002:sink_ready -> APB_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [105:0] syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_003:sink_ready -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [105:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_004:sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                                 // APB_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_valid;                                       // APB_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                               // APB_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [82:0] apb_m0_translator_avalon_universal_master_0_agent_cp_data;                                        // APB_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          apb_m0_translator_avalon_universal_master_0_agent_cp_ready;                                       // addr_router_004:sink_ready -> APB_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [82:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [82:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_006:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [82:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_007:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [82:0] button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_008:sink_ready -> button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [82:0] sw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // sw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_009:sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // hex_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // hex_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // hex_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [82:0] hex_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // hex_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          hex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_010:sink_ready -> hex_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [82:0] motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // motorA_duty_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_011:sink_ready -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [82:0] motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // motorB_duty_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_012:sink_ready -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [82:0] motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // motorA_dir_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_013:sink_ready -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [82:0] motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // motorB_dir_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_014:sink_ready -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // hex_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // hex_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // hex_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [82:0] hex_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // hex_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          hex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_015:sink_ready -> hex_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [82:0] infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_016:sink_ready -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire   [82:0] infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_017:sink_ready -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [82:0] infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_018:sink_ready -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire   [82:0] infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_019:sink_ready -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire   [82:0] infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_020:sink_ready -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_002_src_endofpacket;                                                                  // addr_router_002:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                        // addr_router_002:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                // addr_router_002:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [105:0] addr_router_002_src_data;                                                                         // addr_router_002:src_data -> limiter:cmd_sink_data
	wire    [4:0] addr_router_002_src_channel;                                                                      // addr_router_002:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                        // limiter:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                            // dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                  // addr_router_004:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                        // addr_router_004:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                // addr_router_004:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [82:0] addr_router_004_src_data;                                                                         // addr_router_004:src_data -> limiter_001:cmd_sink_data
	wire   [15:0] addr_router_004_src_channel;                                                                      // addr_router_004:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                        // limiter_001:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                  // limiter_001:rsp_src_endofpacket -> APB_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                        // limiter_001:rsp_src_valid -> APB_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                // limiter_001:rsp_src_startofpacket -> APB_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [82:0] limiter_001_rsp_src_data;                                                                         // limiter_001:rsp_src_data -> APB_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] limiter_001_rsp_src_channel;                                                                      // limiter_001:rsp_src_channel -> APB_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                        // APB_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [87:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                      // sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [4:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                            // burst_adapter_001:source0_endofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                  // burst_adapter_001:source0_valid -> APB_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                          // burst_adapter_001:source0_startofpacket -> APB_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] burst_adapter_001_source0_data;                                                                   // burst_adapter_001:source0_data -> APB_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                  // APB_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [4:0] burst_adapter_001_source0_channel;                                                                // burst_adapter_001:source0_channel -> APB_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [APB:reset, APB_m0_translator:reset, APB_m0_translator_avalon_universal_master_0_agent:reset, APB_s0_translator:reset, APB_s0_translator_avalon_universal_slave_0_agent:reset, APB_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, crosser:in_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, crosser_010:in_reset, crosser_011:in_reset, crosser_012:in_reset, crosser_013:in_reset, crosser_014:in_reset, crosser_015:in_reset, crosser_016:in_reset, crosser_017:in_reset, crosser_018:out_reset, crosser_019:out_reset, crosser_020:out_reset, crosser_021:out_reset, crosser_022:out_reset, crosser_023:out_reset, crosser_024:out_reset, crosser_025:out_reset, crosser_026:out_reset, crosser_027:out_reset, crosser_028:out_reset, crosser_029:out_reset, crosser_030:out_reset, crosser_031:out_reset, crosser_032:out_reset, crosser_033:out_reset, dma:system_reset_n, dma_control_port_slave_translator:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_read_master_translator:reset, dma_read_master_translator_avalon_universal_master_0_agent:reset, dma_write_master_translator:reset, dma_write_master_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_004:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, limiter:reset, limiter_001:reset, nios2cpu:reset_n, nios2cpu_data_master_translator:reset, nios2cpu_data_master_translator_avalon_universal_master_0_agent:reset, nios2cpu_instruction_master_translator:reset, nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2cpu_jtag_debug_module_translator:reset, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_004:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, sdram_ctrl:reset_n, sdram_ctrl_s1_translator:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire          nios2cpu_jtag_debug_module_reset_reset;                                                           // nios2cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [button:reset_n, button_s1_translator:reset, button_s1_translator_avalon_universal_slave_0_agent:reset, button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, crosser_010:out_reset, crosser_011:out_reset, crosser_012:out_reset, crosser_013:out_reset, crosser_014:out_reset, crosser_015:out_reset, crosser_016:out_reset, crosser_017:out_reset, crosser_018:in_reset, crosser_019:in_reset, crosser_020:in_reset, crosser_021:in_reset, crosser_022:in_reset, crosser_023:in_reset, crosser_024:in_reset, crosser_025:in_reset, crosser_026:in_reset, crosser_027:in_reset, crosser_028:in_reset, crosser_029:in_reset, crosser_030:in_reset, crosser_031:in_reset, crosser_032:in_reset, crosser_033:in_reset, hex_0:reset_n, hex_0_s1_translator:reset, hex_0_s1_translator_avalon_universal_slave_0_agent:reset, hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex_1:reset_n, hex_1_s1_translator:reset, hex_1_s1_translator_avalon_universal_slave_0_agent:reset, hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, infra_sensor_0:reset_n, infra_sensor_0_s1_translator:reset, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:reset, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, infra_sensor_1:reset_n, infra_sensor_1_s1_translator:reset, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:reset, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, infra_sensor_2:reset_n, infra_sensor_2_s1_translator:reset, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:reset, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, infra_sensor_3:reset_n, infra_sensor_3_s1_translator:reset, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:reset, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, infra_sensor_4:reset_n, infra_sensor_4_s1_translator:reset, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:reset, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motorA_dir:reset_n, motorA_dir_s1_translator:reset, motorA_dir_s1_translator_avalon_universal_slave_0_agent:reset, motorA_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, motorA_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motorA_duty:reset_n, motorA_duty_s1_translator:reset, motorA_duty_s1_translator_avalon_universal_slave_0_agent:reset, motorA_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, motorA_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motorB_dir:reset_n, motorB_dir_s1_translator:reset, motorB_dir_s1_translator_avalon_universal_slave_0_agent:reset, motorB_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, motorB_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motorB_duty:reset_n, motorB_duty_s1_translator:reset, motorB_duty_s1_translator_avalon_universal_slave_0_agent:reset, motorB_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, motorB_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, sw:reset_n, sw_s1_translator:reset, sw_s1_translator_avalon_universal_slave_0_agent:reset, sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                               // rst_controller_002:reset_out -> [crosser:out_reset, crosser_001:in_reset, id_router_003:reset, rsp_xbar_demux_003:reset, syspll:reset, syspll_pll_slave_translator:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [4:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [4:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [105:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire    [4:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                              // cmd_xbar_demux_001:src4_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                    // cmd_xbar_demux_001:src4_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                            // cmd_xbar_demux_001:src4_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src4_data;                                                                     // cmd_xbar_demux_001:src4_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_001_src4_channel;                                                                  // cmd_xbar_demux_001:src4_channel -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src0_data;                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_001:sink2_data
	wire    [4:0] cmd_xbar_demux_002_src0_channel;                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                    // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                              // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                    // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_002:sink2_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                            // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [105:0] cmd_xbar_demux_002_src1_data;                                                                     // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_002:sink2_data
	wire    [4:0] cmd_xbar_demux_002_src1_channel;                                                                  // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_002:sink2_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                    // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                              // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                    // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                            // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [105:0] cmd_xbar_demux_003_src0_data;                                                                     // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_001:sink3_data
	wire    [4:0] cmd_xbar_demux_003_src0_channel;                                                                  // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                    // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                              // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                    // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_002:sink3_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                            // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	wire  [105:0] cmd_xbar_demux_003_src1_data;                                                                     // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_002:sink3_data
	wire    [4:0] cmd_xbar_demux_003_src1_channel;                                                                  // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_002:sink3_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                    // cmd_xbar_mux_002:sink3_ready -> cmd_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [4:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [4:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                              // rsp_xbar_demux_001:src2_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                    // rsp_xbar_demux_001:src2_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                            // rsp_xbar_demux_001:src2_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src2_data;                                                                     // rsp_xbar_demux_001:src2_data -> rsp_xbar_mux_002:sink0_data
	wire    [4:0] rsp_xbar_demux_001_src2_channel;                                                                  // rsp_xbar_demux_001:src2_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                    // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                              // rsp_xbar_demux_001:src3_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                    // rsp_xbar_demux_001:src3_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                            // rsp_xbar_demux_001:src3_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [105:0] rsp_xbar_demux_001_src3_data;                                                                     // rsp_xbar_demux_001:src3_data -> rsp_xbar_mux_003:sink0_data
	wire    [4:0] rsp_xbar_demux_001_src3_channel;                                                                  // rsp_xbar_demux_001:src3_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_001_src3_ready;                                                                    // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_001:src3_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_002_src2_endofpacket;                                                              // rsp_xbar_demux_002:src2_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_002_src2_valid;                                                                    // rsp_xbar_demux_002:src2_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_002_src2_startofpacket;                                                            // rsp_xbar_demux_002:src2_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src2_data;                                                                     // rsp_xbar_demux_002:src2_data -> rsp_xbar_mux_002:sink1_data
	wire    [4:0] rsp_xbar_demux_002_src2_channel;                                                                  // rsp_xbar_demux_002:src2_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_002_src2_ready;                                                                    // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_002:src2_ready
	wire          rsp_xbar_demux_002_src3_endofpacket;                                                              // rsp_xbar_demux_002:src3_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_002_src3_valid;                                                                    // rsp_xbar_demux_002:src3_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_002_src3_startofpacket;                                                            // rsp_xbar_demux_002:src3_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [105:0] rsp_xbar_demux_002_src3_data;                                                                     // rsp_xbar_demux_002:src3_data -> rsp_xbar_mux_003:sink1_data
	wire    [4:0] rsp_xbar_demux_002_src3_channel;                                                                  // rsp_xbar_demux_002:src3_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_002_src3_ready;                                                                    // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_002:src3_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [105:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [4:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [105:0] addr_router_src_data;                                                                             // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [4:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // nios2cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [105:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [4:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                       // nios2cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [105:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire    [4:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_cmd_src_ready;                                                                            // cmd_xbar_demux_002:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                 // rsp_xbar_mux_002:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                       // rsp_xbar_mux_002:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                               // rsp_xbar_mux_002:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [105:0] rsp_xbar_mux_002_src_data;                                                                        // rsp_xbar_mux_002:src_data -> limiter:rsp_sink_data
	wire    [4:0] rsp_xbar_mux_002_src_channel;                                                                     // rsp_xbar_mux_002:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                       // limiter:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire          addr_router_003_src_endofpacket;                                                                  // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                        // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [105:0] addr_router_003_src_data;                                                                         // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [4:0] addr_router_003_src_channel;                                                                      // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                        // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                 // rsp_xbar_mux_003:src_endofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                       // rsp_xbar_mux_003:src_valid -> dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                               // rsp_xbar_mux_003:src_startofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [105:0] rsp_xbar_mux_003_src_data;                                                                        // rsp_xbar_mux_003:src_data -> dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_003_src_channel;                                                                     // rsp_xbar_mux_003:src_channel -> dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                       // dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_003:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                           // nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [105:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [4:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [105:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> burst_adapter_001:sink0_data
	wire    [4:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                       // burst_adapter_001:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [105:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [4:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          crosser_out_ready;                                                                                // syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [105:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [4:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [105:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [4:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                  // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [82:0] limiter_001_cmd_src_data;                                                                         // limiter_001:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire   [15:0] limiter_001_cmd_src_channel;                                                                      // limiter_001:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                        // cmd_xbar_demux_004:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                 // rsp_xbar_mux_004:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                       // rsp_xbar_mux_004:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                               // rsp_xbar_mux_004:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [82:0] rsp_xbar_mux_004_src_data;                                                                        // rsp_xbar_mux_004:src_data -> limiter_001:rsp_sink_data
	wire   [15:0] rsp_xbar_mux_004_src_channel;                                                                     // rsp_xbar_mux_004:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                       // limiter_001:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	wire          crosser_002_out_ready;                                                                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [82:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [15:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          crosser_003_out_ready;                                                                            // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_003:out_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [82:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [15:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          crosser_004_out_ready;                                                                            // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_004:out_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [82:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [15:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          crosser_005_out_ready;                                                                            // button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_005:out_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [82:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [15:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          crosser_006_out_ready;                                                                            // sw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_006:out_ready
	wire          id_router_009_src_endofpacket;                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [82:0] id_router_009_src_data;                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [15:0] id_router_009_src_channel;                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          crosser_007_out_ready;                                                                            // hex_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_007:out_ready
	wire          id_router_010_src_endofpacket;                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [82:0] id_router_010_src_data;                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [15:0] id_router_010_src_channel;                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          crosser_008_out_ready;                                                                            // motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_008:out_ready
	wire          id_router_011_src_endofpacket;                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [82:0] id_router_011_src_data;                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [15:0] id_router_011_src_channel;                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          crosser_009_out_ready;                                                                            // motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_009:out_ready
	wire          id_router_012_src_endofpacket;                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [82:0] id_router_012_src_data;                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [15:0] id_router_012_src_channel;                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          crosser_010_out_ready;                                                                            // motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_010:out_ready
	wire          id_router_013_src_endofpacket;                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [82:0] id_router_013_src_data;                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [15:0] id_router_013_src_channel;                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          crosser_011_out_ready;                                                                            // motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_011:out_ready
	wire          id_router_014_src_endofpacket;                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [82:0] id_router_014_src_data;                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          crosser_012_out_ready;                                                                            // hex_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_012:out_ready
	wire          id_router_015_src_endofpacket;                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [82:0] id_router_015_src_data;                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          crosser_013_out_ready;                                                                            // infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_013:out_ready
	wire          id_router_016_src_endofpacket;                                                                    // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                          // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                  // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [82:0] id_router_016_src_data;                                                                           // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [15:0] id_router_016_src_channel;                                                                        // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                          // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          crosser_014_out_ready;                                                                            // infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_014:out_ready
	wire          id_router_017_src_endofpacket;                                                                    // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                          // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                  // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire   [82:0] id_router_017_src_data;                                                                           // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [15:0] id_router_017_src_channel;                                                                        // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                          // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          crosser_015_out_ready;                                                                            // infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_015:out_ready
	wire          id_router_018_src_endofpacket;                                                                    // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                          // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                  // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [82:0] id_router_018_src_data;                                                                           // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [15:0] id_router_018_src_channel;                                                                        // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                          // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          crosser_016_out_ready;                                                                            // infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_016:out_ready
	wire          id_router_019_src_endofpacket;                                                                    // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                          // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                  // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire   [82:0] id_router_019_src_data;                                                                           // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [15:0] id_router_019_src_channel;                                                                        // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                          // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          crosser_017_out_ready;                                                                            // infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_017:out_ready
	wire          id_router_020_src_endofpacket;                                                                    // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                          // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                  // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire   [82:0] id_router_020_src_data;                                                                           // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [15:0] id_router_020_src_channel;                                                                        // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                          // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [105:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire    [4:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [87:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [4:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [87:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> width_adapter_001:in_data
	wire    [4:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [105:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire    [4:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          crosser_out_endofpacket;                                                                          // crosser:out_endofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                // crosser:out_valid -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                        // crosser:out_startofpacket -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] crosser_out_data;                                                                                 // crosser:out_data -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] crosser_out_channel;                                                                              // crosser:out_channel -> syspll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> crosser:in_startofpacket
	wire  [105:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> crosser:in_data
	wire    [4:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                    // crosser:in_ready -> cmd_xbar_demux_001:src3_ready
	wire          crosser_001_out_endofpacket;                                                                      // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          crosser_001_out_valid;                                                                            // crosser_001:out_valid -> rsp_xbar_mux_001:sink3_valid
	wire          crosser_001_out_startofpacket;                                                                    // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [105:0] crosser_001_out_data;                                                                             // crosser_001:out_data -> rsp_xbar_mux_001:sink3_data
	wire    [4:0] crosser_001_out_channel;                                                                          // crosser_001:out_channel -> rsp_xbar_mux_001:sink3_channel
	wire          crosser_001_out_ready;                                                                            // rsp_xbar_mux_001:sink3_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [105:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> crosser_001:in_data
	wire    [4:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // crosser_001:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          crosser_002_out_endofpacket;                                                                      // crosser_002:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                            // crosser_002:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                    // crosser_002:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_002_out_data;                                                                             // crosser_002:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_002_out_channel;                                                                          // crosser_002:out_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                              // cmd_xbar_demux_004:src0_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                    // cmd_xbar_demux_004:src0_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                            // cmd_xbar_demux_004:src0_startofpacket -> crosser_002:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src0_data;                                                                     // cmd_xbar_demux_004:src0_data -> crosser_002:in_data
	wire   [15:0] cmd_xbar_demux_004_src0_channel;                                                                  // cmd_xbar_demux_004:src0_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                    // crosser_002:in_ready -> cmd_xbar_demux_004:src0_ready
	wire          crosser_003_out_endofpacket;                                                                      // crosser_003:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_003_out_valid;                                                                            // crosser_003:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_003_out_startofpacket;                                                                    // crosser_003:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_003_out_data;                                                                             // crosser_003:out_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_003_out_channel;                                                                          // crosser_003:out_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                              // cmd_xbar_demux_004:src1_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                    // cmd_xbar_demux_004:src1_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                            // cmd_xbar_demux_004:src1_startofpacket -> crosser_003:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src1_data;                                                                     // cmd_xbar_demux_004:src1_data -> crosser_003:in_data
	wire   [15:0] cmd_xbar_demux_004_src1_channel;                                                                  // cmd_xbar_demux_004:src1_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_004_src1_ready;                                                                    // crosser_003:in_ready -> cmd_xbar_demux_004:src1_ready
	wire          crosser_004_out_endofpacket;                                                                      // crosser_004:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_004_out_valid;                                                                            // crosser_004:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_004_out_startofpacket;                                                                    // crosser_004:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_004_out_data;                                                                             // crosser_004:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_004_out_channel;                                                                          // crosser_004:out_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src2_endofpacket;                                                              // cmd_xbar_demux_004:src2_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_004_src2_valid;                                                                    // cmd_xbar_demux_004:src2_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_004_src2_startofpacket;                                                            // cmd_xbar_demux_004:src2_startofpacket -> crosser_004:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src2_data;                                                                     // cmd_xbar_demux_004:src2_data -> crosser_004:in_data
	wire   [15:0] cmd_xbar_demux_004_src2_channel;                                                                  // cmd_xbar_demux_004:src2_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_004_src2_ready;                                                                    // crosser_004:in_ready -> cmd_xbar_demux_004:src2_ready
	wire          crosser_005_out_endofpacket;                                                                      // crosser_005:out_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_005_out_valid;                                                                            // crosser_005:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_005_out_startofpacket;                                                                    // crosser_005:out_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_005_out_data;                                                                             // crosser_005:out_data -> button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_005_out_channel;                                                                          // crosser_005:out_channel -> button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src3_endofpacket;                                                              // cmd_xbar_demux_004:src3_endofpacket -> crosser_005:in_endofpacket
	wire          cmd_xbar_demux_004_src3_valid;                                                                    // cmd_xbar_demux_004:src3_valid -> crosser_005:in_valid
	wire          cmd_xbar_demux_004_src3_startofpacket;                                                            // cmd_xbar_demux_004:src3_startofpacket -> crosser_005:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src3_data;                                                                     // cmd_xbar_demux_004:src3_data -> crosser_005:in_data
	wire   [15:0] cmd_xbar_demux_004_src3_channel;                                                                  // cmd_xbar_demux_004:src3_channel -> crosser_005:in_channel
	wire          cmd_xbar_demux_004_src3_ready;                                                                    // crosser_005:in_ready -> cmd_xbar_demux_004:src3_ready
	wire          crosser_006_out_endofpacket;                                                                      // crosser_006:out_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_006_out_valid;                                                                            // crosser_006:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_006_out_startofpacket;                                                                    // crosser_006:out_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_006_out_data;                                                                             // crosser_006:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_006_out_channel;                                                                          // crosser_006:out_channel -> sw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src4_endofpacket;                                                              // cmd_xbar_demux_004:src4_endofpacket -> crosser_006:in_endofpacket
	wire          cmd_xbar_demux_004_src4_valid;                                                                    // cmd_xbar_demux_004:src4_valid -> crosser_006:in_valid
	wire          cmd_xbar_demux_004_src4_startofpacket;                                                            // cmd_xbar_demux_004:src4_startofpacket -> crosser_006:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src4_data;                                                                     // cmd_xbar_demux_004:src4_data -> crosser_006:in_data
	wire   [15:0] cmd_xbar_demux_004_src4_channel;                                                                  // cmd_xbar_demux_004:src4_channel -> crosser_006:in_channel
	wire          cmd_xbar_demux_004_src4_ready;                                                                    // crosser_006:in_ready -> cmd_xbar_demux_004:src4_ready
	wire          crosser_007_out_endofpacket;                                                                      // crosser_007:out_endofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_007_out_valid;                                                                            // crosser_007:out_valid -> hex_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_007_out_startofpacket;                                                                    // crosser_007:out_startofpacket -> hex_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_007_out_data;                                                                             // crosser_007:out_data -> hex_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_007_out_channel;                                                                          // crosser_007:out_channel -> hex_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src5_endofpacket;                                                              // cmd_xbar_demux_004:src5_endofpacket -> crosser_007:in_endofpacket
	wire          cmd_xbar_demux_004_src5_valid;                                                                    // cmd_xbar_demux_004:src5_valid -> crosser_007:in_valid
	wire          cmd_xbar_demux_004_src5_startofpacket;                                                            // cmd_xbar_demux_004:src5_startofpacket -> crosser_007:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src5_data;                                                                     // cmd_xbar_demux_004:src5_data -> crosser_007:in_data
	wire   [15:0] cmd_xbar_demux_004_src5_channel;                                                                  // cmd_xbar_demux_004:src5_channel -> crosser_007:in_channel
	wire          cmd_xbar_demux_004_src5_ready;                                                                    // crosser_007:in_ready -> cmd_xbar_demux_004:src5_ready
	wire          crosser_008_out_endofpacket;                                                                      // crosser_008:out_endofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_008_out_valid;                                                                            // crosser_008:out_valid -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_008_out_startofpacket;                                                                    // crosser_008:out_startofpacket -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_008_out_data;                                                                             // crosser_008:out_data -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_008_out_channel;                                                                          // crosser_008:out_channel -> motorA_duty_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src6_endofpacket;                                                              // cmd_xbar_demux_004:src6_endofpacket -> crosser_008:in_endofpacket
	wire          cmd_xbar_demux_004_src6_valid;                                                                    // cmd_xbar_demux_004:src6_valid -> crosser_008:in_valid
	wire          cmd_xbar_demux_004_src6_startofpacket;                                                            // cmd_xbar_demux_004:src6_startofpacket -> crosser_008:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src6_data;                                                                     // cmd_xbar_demux_004:src6_data -> crosser_008:in_data
	wire   [15:0] cmd_xbar_demux_004_src6_channel;                                                                  // cmd_xbar_demux_004:src6_channel -> crosser_008:in_channel
	wire          cmd_xbar_demux_004_src6_ready;                                                                    // crosser_008:in_ready -> cmd_xbar_demux_004:src6_ready
	wire          crosser_009_out_endofpacket;                                                                      // crosser_009:out_endofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_009_out_valid;                                                                            // crosser_009:out_valid -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_009_out_startofpacket;                                                                    // crosser_009:out_startofpacket -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_009_out_data;                                                                             // crosser_009:out_data -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_009_out_channel;                                                                          // crosser_009:out_channel -> motorB_duty_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src7_endofpacket;                                                              // cmd_xbar_demux_004:src7_endofpacket -> crosser_009:in_endofpacket
	wire          cmd_xbar_demux_004_src7_valid;                                                                    // cmd_xbar_demux_004:src7_valid -> crosser_009:in_valid
	wire          cmd_xbar_demux_004_src7_startofpacket;                                                            // cmd_xbar_demux_004:src7_startofpacket -> crosser_009:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src7_data;                                                                     // cmd_xbar_demux_004:src7_data -> crosser_009:in_data
	wire   [15:0] cmd_xbar_demux_004_src7_channel;                                                                  // cmd_xbar_demux_004:src7_channel -> crosser_009:in_channel
	wire          cmd_xbar_demux_004_src7_ready;                                                                    // crosser_009:in_ready -> cmd_xbar_demux_004:src7_ready
	wire          crosser_010_out_endofpacket;                                                                      // crosser_010:out_endofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_010_out_valid;                                                                            // crosser_010:out_valid -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_010_out_startofpacket;                                                                    // crosser_010:out_startofpacket -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_010_out_data;                                                                             // crosser_010:out_data -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_010_out_channel;                                                                          // crosser_010:out_channel -> motorA_dir_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src8_endofpacket;                                                              // cmd_xbar_demux_004:src8_endofpacket -> crosser_010:in_endofpacket
	wire          cmd_xbar_demux_004_src8_valid;                                                                    // cmd_xbar_demux_004:src8_valid -> crosser_010:in_valid
	wire          cmd_xbar_demux_004_src8_startofpacket;                                                            // cmd_xbar_demux_004:src8_startofpacket -> crosser_010:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src8_data;                                                                     // cmd_xbar_demux_004:src8_data -> crosser_010:in_data
	wire   [15:0] cmd_xbar_demux_004_src8_channel;                                                                  // cmd_xbar_demux_004:src8_channel -> crosser_010:in_channel
	wire          cmd_xbar_demux_004_src8_ready;                                                                    // crosser_010:in_ready -> cmd_xbar_demux_004:src8_ready
	wire          crosser_011_out_endofpacket;                                                                      // crosser_011:out_endofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_011_out_valid;                                                                            // crosser_011:out_valid -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_011_out_startofpacket;                                                                    // crosser_011:out_startofpacket -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_011_out_data;                                                                             // crosser_011:out_data -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_011_out_channel;                                                                          // crosser_011:out_channel -> motorB_dir_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src9_endofpacket;                                                              // cmd_xbar_demux_004:src9_endofpacket -> crosser_011:in_endofpacket
	wire          cmd_xbar_demux_004_src9_valid;                                                                    // cmd_xbar_demux_004:src9_valid -> crosser_011:in_valid
	wire          cmd_xbar_demux_004_src9_startofpacket;                                                            // cmd_xbar_demux_004:src9_startofpacket -> crosser_011:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src9_data;                                                                     // cmd_xbar_demux_004:src9_data -> crosser_011:in_data
	wire   [15:0] cmd_xbar_demux_004_src9_channel;                                                                  // cmd_xbar_demux_004:src9_channel -> crosser_011:in_channel
	wire          cmd_xbar_demux_004_src9_ready;                                                                    // crosser_011:in_ready -> cmd_xbar_demux_004:src9_ready
	wire          crosser_012_out_endofpacket;                                                                      // crosser_012:out_endofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_012_out_valid;                                                                            // crosser_012:out_valid -> hex_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_012_out_startofpacket;                                                                    // crosser_012:out_startofpacket -> hex_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_012_out_data;                                                                             // crosser_012:out_data -> hex_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_012_out_channel;                                                                          // crosser_012:out_channel -> hex_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src10_endofpacket;                                                             // cmd_xbar_demux_004:src10_endofpacket -> crosser_012:in_endofpacket
	wire          cmd_xbar_demux_004_src10_valid;                                                                   // cmd_xbar_demux_004:src10_valid -> crosser_012:in_valid
	wire          cmd_xbar_demux_004_src10_startofpacket;                                                           // cmd_xbar_demux_004:src10_startofpacket -> crosser_012:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src10_data;                                                                    // cmd_xbar_demux_004:src10_data -> crosser_012:in_data
	wire   [15:0] cmd_xbar_demux_004_src10_channel;                                                                 // cmd_xbar_demux_004:src10_channel -> crosser_012:in_channel
	wire          cmd_xbar_demux_004_src10_ready;                                                                   // crosser_012:in_ready -> cmd_xbar_demux_004:src10_ready
	wire          crosser_013_out_endofpacket;                                                                      // crosser_013:out_endofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_013_out_valid;                                                                            // crosser_013:out_valid -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_013_out_startofpacket;                                                                    // crosser_013:out_startofpacket -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_013_out_data;                                                                             // crosser_013:out_data -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_013_out_channel;                                                                          // crosser_013:out_channel -> infra_sensor_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src11_endofpacket;                                                             // cmd_xbar_demux_004:src11_endofpacket -> crosser_013:in_endofpacket
	wire          cmd_xbar_demux_004_src11_valid;                                                                   // cmd_xbar_demux_004:src11_valid -> crosser_013:in_valid
	wire          cmd_xbar_demux_004_src11_startofpacket;                                                           // cmd_xbar_demux_004:src11_startofpacket -> crosser_013:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src11_data;                                                                    // cmd_xbar_demux_004:src11_data -> crosser_013:in_data
	wire   [15:0] cmd_xbar_demux_004_src11_channel;                                                                 // cmd_xbar_demux_004:src11_channel -> crosser_013:in_channel
	wire          cmd_xbar_demux_004_src11_ready;                                                                   // crosser_013:in_ready -> cmd_xbar_demux_004:src11_ready
	wire          crosser_014_out_endofpacket;                                                                      // crosser_014:out_endofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_014_out_valid;                                                                            // crosser_014:out_valid -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_014_out_startofpacket;                                                                    // crosser_014:out_startofpacket -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_014_out_data;                                                                             // crosser_014:out_data -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_014_out_channel;                                                                          // crosser_014:out_channel -> infra_sensor_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src12_endofpacket;                                                             // cmd_xbar_demux_004:src12_endofpacket -> crosser_014:in_endofpacket
	wire          cmd_xbar_demux_004_src12_valid;                                                                   // cmd_xbar_demux_004:src12_valid -> crosser_014:in_valid
	wire          cmd_xbar_demux_004_src12_startofpacket;                                                           // cmd_xbar_demux_004:src12_startofpacket -> crosser_014:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src12_data;                                                                    // cmd_xbar_demux_004:src12_data -> crosser_014:in_data
	wire   [15:0] cmd_xbar_demux_004_src12_channel;                                                                 // cmd_xbar_demux_004:src12_channel -> crosser_014:in_channel
	wire          cmd_xbar_demux_004_src12_ready;                                                                   // crosser_014:in_ready -> cmd_xbar_demux_004:src12_ready
	wire          crosser_015_out_endofpacket;                                                                      // crosser_015:out_endofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_015_out_valid;                                                                            // crosser_015:out_valid -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_015_out_startofpacket;                                                                    // crosser_015:out_startofpacket -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_015_out_data;                                                                             // crosser_015:out_data -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_015_out_channel;                                                                          // crosser_015:out_channel -> infra_sensor_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src13_endofpacket;                                                             // cmd_xbar_demux_004:src13_endofpacket -> crosser_015:in_endofpacket
	wire          cmd_xbar_demux_004_src13_valid;                                                                   // cmd_xbar_demux_004:src13_valid -> crosser_015:in_valid
	wire          cmd_xbar_demux_004_src13_startofpacket;                                                           // cmd_xbar_demux_004:src13_startofpacket -> crosser_015:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src13_data;                                                                    // cmd_xbar_demux_004:src13_data -> crosser_015:in_data
	wire   [15:0] cmd_xbar_demux_004_src13_channel;                                                                 // cmd_xbar_demux_004:src13_channel -> crosser_015:in_channel
	wire          cmd_xbar_demux_004_src13_ready;                                                                   // crosser_015:in_ready -> cmd_xbar_demux_004:src13_ready
	wire          crosser_016_out_endofpacket;                                                                      // crosser_016:out_endofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_016_out_valid;                                                                            // crosser_016:out_valid -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_016_out_startofpacket;                                                                    // crosser_016:out_startofpacket -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_016_out_data;                                                                             // crosser_016:out_data -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_016_out_channel;                                                                          // crosser_016:out_channel -> infra_sensor_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src14_endofpacket;                                                             // cmd_xbar_demux_004:src14_endofpacket -> crosser_016:in_endofpacket
	wire          cmd_xbar_demux_004_src14_valid;                                                                   // cmd_xbar_demux_004:src14_valid -> crosser_016:in_valid
	wire          cmd_xbar_demux_004_src14_startofpacket;                                                           // cmd_xbar_demux_004:src14_startofpacket -> crosser_016:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src14_data;                                                                    // cmd_xbar_demux_004:src14_data -> crosser_016:in_data
	wire   [15:0] cmd_xbar_demux_004_src14_channel;                                                                 // cmd_xbar_demux_004:src14_channel -> crosser_016:in_channel
	wire          cmd_xbar_demux_004_src14_ready;                                                                   // crosser_016:in_ready -> cmd_xbar_demux_004:src14_ready
	wire          crosser_017_out_endofpacket;                                                                      // crosser_017:out_endofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_017_out_valid;                                                                            // crosser_017:out_valid -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_017_out_startofpacket;                                                                    // crosser_017:out_startofpacket -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_017_out_data;                                                                             // crosser_017:out_data -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_017_out_channel;                                                                          // crosser_017:out_channel -> infra_sensor_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src15_endofpacket;                                                             // cmd_xbar_demux_004:src15_endofpacket -> crosser_017:in_endofpacket
	wire          cmd_xbar_demux_004_src15_valid;                                                                   // cmd_xbar_demux_004:src15_valid -> crosser_017:in_valid
	wire          cmd_xbar_demux_004_src15_startofpacket;                                                           // cmd_xbar_demux_004:src15_startofpacket -> crosser_017:in_startofpacket
	wire   [82:0] cmd_xbar_demux_004_src15_data;                                                                    // cmd_xbar_demux_004:src15_data -> crosser_017:in_data
	wire   [15:0] cmd_xbar_demux_004_src15_channel;                                                                 // cmd_xbar_demux_004:src15_channel -> crosser_017:in_channel
	wire          cmd_xbar_demux_004_src15_ready;                                                                   // crosser_017:in_ready -> cmd_xbar_demux_004:src15_ready
	wire          crosser_018_out_endofpacket;                                                                      // crosser_018:out_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          crosser_018_out_valid;                                                                            // crosser_018:out_valid -> rsp_xbar_mux_004:sink0_valid
	wire          crosser_018_out_startofpacket;                                                                    // crosser_018:out_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire   [82:0] crosser_018_out_data;                                                                             // crosser_018:out_data -> rsp_xbar_mux_004:sink0_data
	wire   [15:0] crosser_018_out_channel;                                                                          // crosser_018:out_channel -> rsp_xbar_mux_004:sink0_channel
	wire          crosser_018_out_ready;                                                                            // rsp_xbar_mux_004:sink0_ready -> crosser_018:out_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> crosser_018:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> crosser_018:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> crosser_018:in_startofpacket
	wire   [82:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> crosser_018:in_data
	wire   [15:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> crosser_018:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // crosser_018:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          crosser_019_out_endofpacket;                                                                      // crosser_019:out_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          crosser_019_out_valid;                                                                            // crosser_019:out_valid -> rsp_xbar_mux_004:sink1_valid
	wire          crosser_019_out_startofpacket;                                                                    // crosser_019:out_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire   [82:0] crosser_019_out_data;                                                                             // crosser_019:out_data -> rsp_xbar_mux_004:sink1_data
	wire   [15:0] crosser_019_out_channel;                                                                          // crosser_019:out_channel -> rsp_xbar_mux_004:sink1_channel
	wire          crosser_019_out_ready;                                                                            // rsp_xbar_mux_004:sink1_ready -> crosser_019:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> crosser_019:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> crosser_019:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> crosser_019:in_startofpacket
	wire   [82:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> crosser_019:in_data
	wire   [15:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> crosser_019:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // crosser_019:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          crosser_020_out_endofpacket;                                                                      // crosser_020:out_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire          crosser_020_out_valid;                                                                            // crosser_020:out_valid -> rsp_xbar_mux_004:sink2_valid
	wire          crosser_020_out_startofpacket;                                                                    // crosser_020:out_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire   [82:0] crosser_020_out_data;                                                                             // crosser_020:out_data -> rsp_xbar_mux_004:sink2_data
	wire   [15:0] crosser_020_out_channel;                                                                          // crosser_020:out_channel -> rsp_xbar_mux_004:sink2_channel
	wire          crosser_020_out_ready;                                                                            // rsp_xbar_mux_004:sink2_ready -> crosser_020:out_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> crosser_020:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> crosser_020:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> crosser_020:in_startofpacket
	wire   [82:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> crosser_020:in_data
	wire   [15:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> crosser_020:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // crosser_020:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          crosser_021_out_endofpacket;                                                                      // crosser_021:out_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	wire          crosser_021_out_valid;                                                                            // crosser_021:out_valid -> rsp_xbar_mux_004:sink3_valid
	wire          crosser_021_out_startofpacket;                                                                    // crosser_021:out_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	wire   [82:0] crosser_021_out_data;                                                                             // crosser_021:out_data -> rsp_xbar_mux_004:sink3_data
	wire   [15:0] crosser_021_out_channel;                                                                          // crosser_021:out_channel -> rsp_xbar_mux_004:sink3_channel
	wire          crosser_021_out_ready;                                                                            // rsp_xbar_mux_004:sink3_ready -> crosser_021:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> crosser_021:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> crosser_021:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> crosser_021:in_startofpacket
	wire   [82:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> crosser_021:in_data
	wire   [15:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> crosser_021:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // crosser_021:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_022_out_endofpacket;                                                                      // crosser_022:out_endofpacket -> rsp_xbar_mux_004:sink4_endofpacket
	wire          crosser_022_out_valid;                                                                            // crosser_022:out_valid -> rsp_xbar_mux_004:sink4_valid
	wire          crosser_022_out_startofpacket;                                                                    // crosser_022:out_startofpacket -> rsp_xbar_mux_004:sink4_startofpacket
	wire   [82:0] crosser_022_out_data;                                                                             // crosser_022:out_data -> rsp_xbar_mux_004:sink4_data
	wire   [15:0] crosser_022_out_channel;                                                                          // crosser_022:out_channel -> rsp_xbar_mux_004:sink4_channel
	wire          crosser_022_out_ready;                                                                            // rsp_xbar_mux_004:sink4_ready -> crosser_022:out_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                              // rsp_xbar_demux_009:src0_endofpacket -> crosser_022:in_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                    // rsp_xbar_demux_009:src0_valid -> crosser_022:in_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                            // rsp_xbar_demux_009:src0_startofpacket -> crosser_022:in_startofpacket
	wire   [82:0] rsp_xbar_demux_009_src0_data;                                                                     // rsp_xbar_demux_009:src0_data -> crosser_022:in_data
	wire   [15:0] rsp_xbar_demux_009_src0_channel;                                                                  // rsp_xbar_demux_009:src0_channel -> crosser_022:in_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                    // crosser_022:in_ready -> rsp_xbar_demux_009:src0_ready
	wire          crosser_023_out_endofpacket;                                                                      // crosser_023:out_endofpacket -> rsp_xbar_mux_004:sink5_endofpacket
	wire          crosser_023_out_valid;                                                                            // crosser_023:out_valid -> rsp_xbar_mux_004:sink5_valid
	wire          crosser_023_out_startofpacket;                                                                    // crosser_023:out_startofpacket -> rsp_xbar_mux_004:sink5_startofpacket
	wire   [82:0] crosser_023_out_data;                                                                             // crosser_023:out_data -> rsp_xbar_mux_004:sink5_data
	wire   [15:0] crosser_023_out_channel;                                                                          // crosser_023:out_channel -> rsp_xbar_mux_004:sink5_channel
	wire          crosser_023_out_ready;                                                                            // rsp_xbar_mux_004:sink5_ready -> crosser_023:out_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                              // rsp_xbar_demux_010:src0_endofpacket -> crosser_023:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                    // rsp_xbar_demux_010:src0_valid -> crosser_023:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                            // rsp_xbar_demux_010:src0_startofpacket -> crosser_023:in_startofpacket
	wire   [82:0] rsp_xbar_demux_010_src0_data;                                                                     // rsp_xbar_demux_010:src0_data -> crosser_023:in_data
	wire   [15:0] rsp_xbar_demux_010_src0_channel;                                                                  // rsp_xbar_demux_010:src0_channel -> crosser_023:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                    // crosser_023:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          crosser_024_out_endofpacket;                                                                      // crosser_024:out_endofpacket -> rsp_xbar_mux_004:sink6_endofpacket
	wire          crosser_024_out_valid;                                                                            // crosser_024:out_valid -> rsp_xbar_mux_004:sink6_valid
	wire          crosser_024_out_startofpacket;                                                                    // crosser_024:out_startofpacket -> rsp_xbar_mux_004:sink6_startofpacket
	wire   [82:0] crosser_024_out_data;                                                                             // crosser_024:out_data -> rsp_xbar_mux_004:sink6_data
	wire   [15:0] crosser_024_out_channel;                                                                          // crosser_024:out_channel -> rsp_xbar_mux_004:sink6_channel
	wire          crosser_024_out_ready;                                                                            // rsp_xbar_mux_004:sink6_ready -> crosser_024:out_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                              // rsp_xbar_demux_011:src0_endofpacket -> crosser_024:in_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                    // rsp_xbar_demux_011:src0_valid -> crosser_024:in_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                            // rsp_xbar_demux_011:src0_startofpacket -> crosser_024:in_startofpacket
	wire   [82:0] rsp_xbar_demux_011_src0_data;                                                                     // rsp_xbar_demux_011:src0_data -> crosser_024:in_data
	wire   [15:0] rsp_xbar_demux_011_src0_channel;                                                                  // rsp_xbar_demux_011:src0_channel -> crosser_024:in_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                    // crosser_024:in_ready -> rsp_xbar_demux_011:src0_ready
	wire          crosser_025_out_endofpacket;                                                                      // crosser_025:out_endofpacket -> rsp_xbar_mux_004:sink7_endofpacket
	wire          crosser_025_out_valid;                                                                            // crosser_025:out_valid -> rsp_xbar_mux_004:sink7_valid
	wire          crosser_025_out_startofpacket;                                                                    // crosser_025:out_startofpacket -> rsp_xbar_mux_004:sink7_startofpacket
	wire   [82:0] crosser_025_out_data;                                                                             // crosser_025:out_data -> rsp_xbar_mux_004:sink7_data
	wire   [15:0] crosser_025_out_channel;                                                                          // crosser_025:out_channel -> rsp_xbar_mux_004:sink7_channel
	wire          crosser_025_out_ready;                                                                            // rsp_xbar_mux_004:sink7_ready -> crosser_025:out_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                              // rsp_xbar_demux_012:src0_endofpacket -> crosser_025:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                    // rsp_xbar_demux_012:src0_valid -> crosser_025:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                            // rsp_xbar_demux_012:src0_startofpacket -> crosser_025:in_startofpacket
	wire   [82:0] rsp_xbar_demux_012_src0_data;                                                                     // rsp_xbar_demux_012:src0_data -> crosser_025:in_data
	wire   [15:0] rsp_xbar_demux_012_src0_channel;                                                                  // rsp_xbar_demux_012:src0_channel -> crosser_025:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                    // crosser_025:in_ready -> rsp_xbar_demux_012:src0_ready
	wire          crosser_026_out_endofpacket;                                                                      // crosser_026:out_endofpacket -> rsp_xbar_mux_004:sink8_endofpacket
	wire          crosser_026_out_valid;                                                                            // crosser_026:out_valid -> rsp_xbar_mux_004:sink8_valid
	wire          crosser_026_out_startofpacket;                                                                    // crosser_026:out_startofpacket -> rsp_xbar_mux_004:sink8_startofpacket
	wire   [82:0] crosser_026_out_data;                                                                             // crosser_026:out_data -> rsp_xbar_mux_004:sink8_data
	wire   [15:0] crosser_026_out_channel;                                                                          // crosser_026:out_channel -> rsp_xbar_mux_004:sink8_channel
	wire          crosser_026_out_ready;                                                                            // rsp_xbar_mux_004:sink8_ready -> crosser_026:out_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                              // rsp_xbar_demux_013:src0_endofpacket -> crosser_026:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                    // rsp_xbar_demux_013:src0_valid -> crosser_026:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                            // rsp_xbar_demux_013:src0_startofpacket -> crosser_026:in_startofpacket
	wire   [82:0] rsp_xbar_demux_013_src0_data;                                                                     // rsp_xbar_demux_013:src0_data -> crosser_026:in_data
	wire   [15:0] rsp_xbar_demux_013_src0_channel;                                                                  // rsp_xbar_demux_013:src0_channel -> crosser_026:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                    // crosser_026:in_ready -> rsp_xbar_demux_013:src0_ready
	wire          crosser_027_out_endofpacket;                                                                      // crosser_027:out_endofpacket -> rsp_xbar_mux_004:sink9_endofpacket
	wire          crosser_027_out_valid;                                                                            // crosser_027:out_valid -> rsp_xbar_mux_004:sink9_valid
	wire          crosser_027_out_startofpacket;                                                                    // crosser_027:out_startofpacket -> rsp_xbar_mux_004:sink9_startofpacket
	wire   [82:0] crosser_027_out_data;                                                                             // crosser_027:out_data -> rsp_xbar_mux_004:sink9_data
	wire   [15:0] crosser_027_out_channel;                                                                          // crosser_027:out_channel -> rsp_xbar_mux_004:sink9_channel
	wire          crosser_027_out_ready;                                                                            // rsp_xbar_mux_004:sink9_ready -> crosser_027:out_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                              // rsp_xbar_demux_014:src0_endofpacket -> crosser_027:in_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                    // rsp_xbar_demux_014:src0_valid -> crosser_027:in_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                            // rsp_xbar_demux_014:src0_startofpacket -> crosser_027:in_startofpacket
	wire   [82:0] rsp_xbar_demux_014_src0_data;                                                                     // rsp_xbar_demux_014:src0_data -> crosser_027:in_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                  // rsp_xbar_demux_014:src0_channel -> crosser_027:in_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                    // crosser_027:in_ready -> rsp_xbar_demux_014:src0_ready
	wire          crosser_028_out_endofpacket;                                                                      // crosser_028:out_endofpacket -> rsp_xbar_mux_004:sink10_endofpacket
	wire          crosser_028_out_valid;                                                                            // crosser_028:out_valid -> rsp_xbar_mux_004:sink10_valid
	wire          crosser_028_out_startofpacket;                                                                    // crosser_028:out_startofpacket -> rsp_xbar_mux_004:sink10_startofpacket
	wire   [82:0] crosser_028_out_data;                                                                             // crosser_028:out_data -> rsp_xbar_mux_004:sink10_data
	wire   [15:0] crosser_028_out_channel;                                                                          // crosser_028:out_channel -> rsp_xbar_mux_004:sink10_channel
	wire          crosser_028_out_ready;                                                                            // rsp_xbar_mux_004:sink10_ready -> crosser_028:out_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                              // rsp_xbar_demux_015:src0_endofpacket -> crosser_028:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                    // rsp_xbar_demux_015:src0_valid -> crosser_028:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                            // rsp_xbar_demux_015:src0_startofpacket -> crosser_028:in_startofpacket
	wire   [82:0] rsp_xbar_demux_015_src0_data;                                                                     // rsp_xbar_demux_015:src0_data -> crosser_028:in_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                  // rsp_xbar_demux_015:src0_channel -> crosser_028:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                    // crosser_028:in_ready -> rsp_xbar_demux_015:src0_ready
	wire          crosser_029_out_endofpacket;                                                                      // crosser_029:out_endofpacket -> rsp_xbar_mux_004:sink11_endofpacket
	wire          crosser_029_out_valid;                                                                            // crosser_029:out_valid -> rsp_xbar_mux_004:sink11_valid
	wire          crosser_029_out_startofpacket;                                                                    // crosser_029:out_startofpacket -> rsp_xbar_mux_004:sink11_startofpacket
	wire   [82:0] crosser_029_out_data;                                                                             // crosser_029:out_data -> rsp_xbar_mux_004:sink11_data
	wire   [15:0] crosser_029_out_channel;                                                                          // crosser_029:out_channel -> rsp_xbar_mux_004:sink11_channel
	wire          crosser_029_out_ready;                                                                            // rsp_xbar_mux_004:sink11_ready -> crosser_029:out_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                              // rsp_xbar_demux_016:src0_endofpacket -> crosser_029:in_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                    // rsp_xbar_demux_016:src0_valid -> crosser_029:in_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                            // rsp_xbar_demux_016:src0_startofpacket -> crosser_029:in_startofpacket
	wire   [82:0] rsp_xbar_demux_016_src0_data;                                                                     // rsp_xbar_demux_016:src0_data -> crosser_029:in_data
	wire   [15:0] rsp_xbar_demux_016_src0_channel;                                                                  // rsp_xbar_demux_016:src0_channel -> crosser_029:in_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                    // crosser_029:in_ready -> rsp_xbar_demux_016:src0_ready
	wire          crosser_030_out_endofpacket;                                                                      // crosser_030:out_endofpacket -> rsp_xbar_mux_004:sink12_endofpacket
	wire          crosser_030_out_valid;                                                                            // crosser_030:out_valid -> rsp_xbar_mux_004:sink12_valid
	wire          crosser_030_out_startofpacket;                                                                    // crosser_030:out_startofpacket -> rsp_xbar_mux_004:sink12_startofpacket
	wire   [82:0] crosser_030_out_data;                                                                             // crosser_030:out_data -> rsp_xbar_mux_004:sink12_data
	wire   [15:0] crosser_030_out_channel;                                                                          // crosser_030:out_channel -> rsp_xbar_mux_004:sink12_channel
	wire          crosser_030_out_ready;                                                                            // rsp_xbar_mux_004:sink12_ready -> crosser_030:out_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                              // rsp_xbar_demux_017:src0_endofpacket -> crosser_030:in_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                    // rsp_xbar_demux_017:src0_valid -> crosser_030:in_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                            // rsp_xbar_demux_017:src0_startofpacket -> crosser_030:in_startofpacket
	wire   [82:0] rsp_xbar_demux_017_src0_data;                                                                     // rsp_xbar_demux_017:src0_data -> crosser_030:in_data
	wire   [15:0] rsp_xbar_demux_017_src0_channel;                                                                  // rsp_xbar_demux_017:src0_channel -> crosser_030:in_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                    // crosser_030:in_ready -> rsp_xbar_demux_017:src0_ready
	wire          crosser_031_out_endofpacket;                                                                      // crosser_031:out_endofpacket -> rsp_xbar_mux_004:sink13_endofpacket
	wire          crosser_031_out_valid;                                                                            // crosser_031:out_valid -> rsp_xbar_mux_004:sink13_valid
	wire          crosser_031_out_startofpacket;                                                                    // crosser_031:out_startofpacket -> rsp_xbar_mux_004:sink13_startofpacket
	wire   [82:0] crosser_031_out_data;                                                                             // crosser_031:out_data -> rsp_xbar_mux_004:sink13_data
	wire   [15:0] crosser_031_out_channel;                                                                          // crosser_031:out_channel -> rsp_xbar_mux_004:sink13_channel
	wire          crosser_031_out_ready;                                                                            // rsp_xbar_mux_004:sink13_ready -> crosser_031:out_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                              // rsp_xbar_demux_018:src0_endofpacket -> crosser_031:in_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                    // rsp_xbar_demux_018:src0_valid -> crosser_031:in_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                            // rsp_xbar_demux_018:src0_startofpacket -> crosser_031:in_startofpacket
	wire   [82:0] rsp_xbar_demux_018_src0_data;                                                                     // rsp_xbar_demux_018:src0_data -> crosser_031:in_data
	wire   [15:0] rsp_xbar_demux_018_src0_channel;                                                                  // rsp_xbar_demux_018:src0_channel -> crosser_031:in_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                    // crosser_031:in_ready -> rsp_xbar_demux_018:src0_ready
	wire          crosser_032_out_endofpacket;                                                                      // crosser_032:out_endofpacket -> rsp_xbar_mux_004:sink14_endofpacket
	wire          crosser_032_out_valid;                                                                            // crosser_032:out_valid -> rsp_xbar_mux_004:sink14_valid
	wire          crosser_032_out_startofpacket;                                                                    // crosser_032:out_startofpacket -> rsp_xbar_mux_004:sink14_startofpacket
	wire   [82:0] crosser_032_out_data;                                                                             // crosser_032:out_data -> rsp_xbar_mux_004:sink14_data
	wire   [15:0] crosser_032_out_channel;                                                                          // crosser_032:out_channel -> rsp_xbar_mux_004:sink14_channel
	wire          crosser_032_out_ready;                                                                            // rsp_xbar_mux_004:sink14_ready -> crosser_032:out_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                              // rsp_xbar_demux_019:src0_endofpacket -> crosser_032:in_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                    // rsp_xbar_demux_019:src0_valid -> crosser_032:in_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                            // rsp_xbar_demux_019:src0_startofpacket -> crosser_032:in_startofpacket
	wire   [82:0] rsp_xbar_demux_019_src0_data;                                                                     // rsp_xbar_demux_019:src0_data -> crosser_032:in_data
	wire   [15:0] rsp_xbar_demux_019_src0_channel;                                                                  // rsp_xbar_demux_019:src0_channel -> crosser_032:in_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                    // crosser_032:in_ready -> rsp_xbar_demux_019:src0_ready
	wire          crosser_033_out_endofpacket;                                                                      // crosser_033:out_endofpacket -> rsp_xbar_mux_004:sink15_endofpacket
	wire          crosser_033_out_valid;                                                                            // crosser_033:out_valid -> rsp_xbar_mux_004:sink15_valid
	wire          crosser_033_out_startofpacket;                                                                    // crosser_033:out_startofpacket -> rsp_xbar_mux_004:sink15_startofpacket
	wire   [82:0] crosser_033_out_data;                                                                             // crosser_033:out_data -> rsp_xbar_mux_004:sink15_data
	wire   [15:0] crosser_033_out_channel;                                                                          // crosser_033:out_channel -> rsp_xbar_mux_004:sink15_channel
	wire          crosser_033_out_ready;                                                                            // rsp_xbar_mux_004:sink15_ready -> crosser_033:out_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                              // rsp_xbar_demux_020:src0_endofpacket -> crosser_033:in_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                    // rsp_xbar_demux_020:src0_valid -> crosser_033:in_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                            // rsp_xbar_demux_020:src0_startofpacket -> crosser_033:in_startofpacket
	wire   [82:0] rsp_xbar_demux_020_src0_data;                                                                     // rsp_xbar_demux_020:src0_data -> crosser_033:in_data
	wire   [15:0] rsp_xbar_demux_020_src0_channel;                                                                  // rsp_xbar_demux_020:src0_channel -> crosser_033:in_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                    // crosser_033:in_ready -> rsp_xbar_demux_020:src0_ready
	wire    [4:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire   [15:0] limiter_001_cmd_valid_data;                                                                       // limiter_001:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                         // dma:dma_ctl_irq -> irq_mapper:receiver0_irq
	wire   [31:0] nios2cpu_d_irq_irq;                                                                               // irq_mapper:sender_irq -> nios2cpu:d_irq
	wire          irq_mapper_receiver1_irq;                                                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                    // jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                // timer:irq -> irq_synchronizer_001:receiver_irq

	DE0Qsys_nios2cpu nios2cpu (
		.clk                                   (syspll_c0_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                       //                   reset_n.reset_n
		.d_address                             (nios2cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2cpu_data_master_read),                                             //                          .read
		.d_readdata                            (nios2cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2cpu_data_master_write),                                            //                          .write
		.d_writedata                           (nios2cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                       // custom_instruction_master.readra
	);

	DE0Qsys_jtag_uart jtag_uart (
		.clk            (syspll_c2_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                                           //               irq.irq
	);

	DE0Qsys_syspll syspll (
		.clk       (clk_50m_clk),                                               //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),                        // inclk_interface_reset.reset
		.read      (syspll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (syspll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (syspll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (syspll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (syspll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (syspll_c0_clk),                                             //                    c0.clk
		.c1        (dram_clk_clk),                                              //                    c1.clk
		.c2        (syspll_c2_clk),                                             //                    c2.clk
		.areset    (areset_export),                                             //        areset_conduit.export
		.locked    (locked_export),                                             //        locked_conduit.export
		.phasedone (phasedone_export)                                           //     phasedone_conduit.export
	);

	DE0Qsys_sdram_ctrl sdram_ctrl (
		.clk            (syspll_c0_clk),                                              //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                            // reset.reset_n
		.az_addr        (sdram_ctrl_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_ctrl_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wires_addr),                                           //  wire.export
		.zs_ba          (sdram_wires_ba),                                             //      .export
		.zs_cas_n       (sdram_wires_cas_n),                                          //      .export
		.zs_cke         (sdram_wires_cke),                                            //      .export
		.zs_cs_n        (sdram_wires_cs_n),                                           //      .export
		.zs_dq          (sdram_wires_dq),                                             //      .export
		.zs_dqm         (sdram_wires_dqm),                                            //      .export
		.zs_ras_n       (sdram_wires_ras_n),                                          //      .export
		.zs_we_n        (sdram_wires_we_n)                                            //      .export
	);

	DE0Qsys_led led (
		.clk        (syspll_c2_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                        // external_connection.export
	);

	DE0Qsys_dma dma (
		.clk                (syspll_c0_clk),                                                    //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                  //              reset.reset_n
		.dma_ctl_address    (dma_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver0_irq),                                         //                irq.irq
		.read_address       (dma_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_read_master_waitrequest),                                      //                   .waitrequest
		.read_burstcount    (dma_read_master_burstcount),                                       //                   .burstcount
		.write_address      (dma_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_write_master_byteenable),                                      //                   .byteenable
		.write_burstcount   (dma_write_master_burstcount)                                       //                   .burstcount
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) apb (
		.clk              (syspll_c0_clk),                                       //   clk.clk
		.reset            (rst_controller_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (apb_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (apb_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (apb_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (apb_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (apb_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (apb_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (apb_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (apb_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (apb_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (apb_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (apb_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (apb_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (apb_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (apb_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (apb_m0_writedata),                                    //      .writedata
		.m0_address       (apb_m0_address),                                      //      .address
		.m0_write         (apb_m0_write),                                        //      .write
		.m0_read          (apb_m0_read),                                         //      .read
		.m0_byteenable    (apb_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (apb_m0_debugaccess)                                   //      .debugaccess
	);

	DE0Qsys_timer timer (
		.clk        (syspll_c2_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                   //   irq.irq
	);

	DE0Qsys_button button (
		.clk        (syspll_c2_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (button_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (button_export)                                        // external_connection.export
	);

	DE0Qsys_sw sw (
		.clk        (syspll_c2_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (sw_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sw_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sw_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sw_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sw_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (sw_export)                                        // external_connection.export
	);

	DE0Qsys_hex_0 hex_0 (
		.clk        (syspll_c2_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address    (hex_0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex_0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex_0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex_0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex_0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex_0_export)                                        // external_connection.export
	);

	DE0Qsys_hex_0 motora_duty (
		.clk        (syspll_c2_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (motora_duty_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~motora_duty_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (motora_duty_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (motora_duty_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (motora_duty_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (motora_duty_export)                                        // external_connection.export
	);

	DE0Qsys_hex_0 motorb_duty (
		.clk        (syspll_c2_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (motorb_duty_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~motorb_duty_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (motorb_duty_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (motorb_duty_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (motorb_duty_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (motorb_duty_export)                                        // external_connection.export
	);

	DE0Qsys_motorA_dir motora_dir (
		.clk        (syspll_c2_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (motora_dir_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~motora_dir_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (motora_dir_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (motora_dir_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (motora_dir_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (motora_dir_export)                                        // external_connection.export
	);

	DE0Qsys_motorA_dir motorb_dir (
		.clk        (syspll_c2_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (motorb_dir_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~motorb_dir_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (motorb_dir_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (motorb_dir_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (motorb_dir_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (motorb_dir_export)                                        // external_connection.export
	);

	DE0Qsys_hex_0 hex_1 (
		.clk        (syspll_c2_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address    (hex_1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex_1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex_1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex_1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex_1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex_1_export)                                        // external_connection.export
	);

	DE0Qsys_infra_sensor_0 infra_sensor_0 (
		.clk      (syspll_c2_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address  (infra_sensor_0_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (infra_sensor_0_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (infra_sensor_0_export)                                      // external_connection.export
	);

	DE0Qsys_infra_sensor_0 infra_sensor_1 (
		.clk      (syspll_c2_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address  (infra_sensor_1_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (infra_sensor_1_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (infra_sensor_1_export)                                      // external_connection.export
	);

	DE0Qsys_infra_sensor_0 infra_sensor_2 (
		.clk      (syspll_c2_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address  (infra_sensor_2_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (infra_sensor_2_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (infra_sensor_2_export)                                      // external_connection.export
	);

	DE0Qsys_infra_sensor_0 infra_sensor_3 (
		.clk      (syspll_c2_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address  (infra_sensor_3_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (infra_sensor_3_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (infra_sensor_3_export)                                      // external_connection.export
	);

	DE0Qsys_infra_sensor_0 infra_sensor_4 (
		.clk      (syspll_c2_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address  (infra_sensor_4_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (infra_sensor_4_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (infra_sensor_4_export)                                      // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2cpu_instruction_master_translator (
		.clk                      (syspll_c0_clk),                                                                  //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address              (nios2cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_byteenable            (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2cpu_data_master_translator (
		.clk                      (syspll_c0_clk),                                                           //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address              (nios2cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2cpu_data_master_read),                                               //                          .read
		.av_readdata              (nios2cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2cpu_data_master_write),                                              //                          .write
		.av_writedata             (nios2cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (8),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_read_master_translator (
		.clk                      (syspll_c0_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_read_master_burstcount),                                         //                          .burstcount
		.av_chipselect            (dma_read_master_chipselect),                                         //                          .chipselect
		.av_read                  (~dma_read_master_read),                                              //                          .read
		.av_readdata              (dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_write                 (1'b0),                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (8),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_write_master_translator (
		.clk                      (syspll_c0_clk),                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address              (dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_write_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (dma_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_write_master_write),                                             //                          .write
		.av_writedata             (dma_write_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                                //               (terminated)
		.av_begintransfer         (1'b0),                                                                //               (terminated)
		.av_read                  (1'b0),                                                                //               (terminated)
		.av_readdata              (),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                //               (terminated)
		.av_debugaccess           (1'b0),                                                                //               (terminated)
		.uav_clken                (),                                                                    //               (terminated)
		.av_clken                 (1'b1),                                                                //               (terminated)
		.uav_response             (2'b00),                                                               //               (terminated)
		.av_response              (),                                                                    //               (terminated)
		.uav_writeresponserequest (),                                                                    //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                //               (terminated)
		.av_writeresponsevalid    ()                                                                     //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2cpu_jtag_debug_module_translator (
		.clk                      (syspll_c0_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_ctrl_s1_translator (
		.clk                      (syspll_c0_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_ctrl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_ctrl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_ctrl_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_ctrl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_ctrl_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_ctrl_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_ctrl_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_ctrl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) apb_s0_translator (
		.clk                      (syspll_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (apb_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (apb_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (apb_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (apb_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (apb_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (apb_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (apb_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (apb_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (apb_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (apb_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (apb_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (apb_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_chipselect            (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) syspll_pll_slave_translator (
		.clk                      (clk_50m_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address              (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (syspll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (syspll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (syspll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (syspll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (syspll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_chipselect            (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (26),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_control_port_slave_translator (
		.clk                      (syspll_c0_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                  //              (terminated)
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) apb_m0_translator (
		.clk                      (syspll_c0_clk),                                             //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                            //                     reset.reset
		.uav_address              (apb_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (apb_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (apb_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (apb_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (apb_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (apb_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (apb_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (apb_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (apb_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (apb_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (apb_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (apb_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (apb_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (apb_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (apb_m0_byteenable),                                         //                          .byteenable
		.av_read                  (apb_m0_read),                                               //                          .read
		.av_readdata              (apb_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (apb_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (apb_m0_write),                                              //                          .write
		.av_writedata             (apb_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (apb_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                      //               (terminated)
		.av_lock                  (1'b0),                                                      //               (terminated)
		.uav_clken                (),                                                          //               (terminated)
		.av_clken                 (1'b1),                                                      //               (terminated)
		.uav_response             (2'b00),                                                     //               (terminated)
		.av_response              (),                                                          //               (terminated)
		.uav_writeresponserequest (),                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (syspll_c2_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (syspll_c2_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (syspll_c2_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_s1_translator (
		.clk                      (syspll_c2_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (button_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (button_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (button_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_s1_translator (
		.clk                      (syspll_c2_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                               //                    reset.reset
		.uav_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sw_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sw_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sw_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                 //              (terminated)
		.av_begintransfer         (),                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                 //              (terminated)
		.av_burstcount            (),                                                                 //              (terminated)
		.av_byteenable            (),                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                             //              (terminated)
		.av_writebyteenable       (),                                                                 //              (terminated)
		.av_lock                  (),                                                                 //              (terminated)
		.av_clken                 (),                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                             //              (terminated)
		.av_debugaccess           (),                                                                 //              (terminated)
		.av_outputenable          (),                                                                 //              (terminated)
		.uav_response             (),                                                                 //              (terminated)
		.av_response              (2'b00),                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex_0_s1_translator (
		.clk                      (syspll_c2_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) motora_duty_s1_translator (
		.clk                      (syspll_c2_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (motora_duty_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (motora_duty_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (motora_duty_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (motora_duty_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (motora_duty_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) motorb_duty_s1_translator (
		.clk                      (syspll_c2_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (motorb_duty_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (motorb_duty_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (motorb_duty_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (motorb_duty_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (motorb_duty_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) motora_dir_s1_translator (
		.clk                      (syspll_c2_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (motora_dir_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (motora_dir_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (motora_dir_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (motora_dir_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (motora_dir_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) motorb_dir_s1_translator (
		.clk                      (syspll_c2_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (motorb_dir_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (motorb_dir_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (motorb_dir_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (motorb_dir_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (motorb_dir_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex_1_s1_translator (
		.clk                      (syspll_c2_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) infra_sensor_0_s1_translator (
		.clk                      (syspll_c2_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (infra_sensor_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (infra_sensor_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                             //              (terminated)
		.av_read                  (),                                                                             //              (terminated)
		.av_writedata             (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) infra_sensor_1_s1_translator (
		.clk                      (syspll_c2_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (infra_sensor_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (infra_sensor_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                             //              (terminated)
		.av_read                  (),                                                                             //              (terminated)
		.av_writedata             (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) infra_sensor_2_s1_translator (
		.clk                      (syspll_c2_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (infra_sensor_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (infra_sensor_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                             //              (terminated)
		.av_read                  (),                                                                             //              (terminated)
		.av_writedata             (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) infra_sensor_3_s1_translator (
		.clk                      (syspll_c2_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (infra_sensor_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (infra_sensor_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                             //              (terminated)
		.av_read                  (),                                                                             //              (terminated)
		.av_writedata             (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) infra_sensor_4_s1_translator (
		.clk                      (syspll_c2_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (infra_sensor_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (infra_sensor_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                             //              (terminated)
		.av_read                  (),                                                                             //              (terminated)
		.av_writedata             (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                           //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address              (nios2cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                   //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                  //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                    //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (nios2cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                       //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                        //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                     //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                       //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                               //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                       //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (96),
		.PKT_THREAD_ID_L           (96),
		.PKT_CACHE_H               (103),
		.PKT_CACHE_L               (100),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address              (dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_003_src_valid),                                                   //        rp.valid
		.rp_data                 (rsp_xbar_mux_003_src_data),                                                    //          .data
		.rp_channel              (rsp_xbar_mux_003_src_channel),                                                 //          .channel
		.rp_startofpacket        (rsp_xbar_mux_003_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_003_src_endofpacket),                                             //          .endofpacket
		.rp_ready                (rsp_xbar_mux_003_src_ready),                                                   //          .ready
		.av_response             (),                                                                             // (terminated)
		.av_writeresponserequest (1'b0),                                                                         // (terminated)
		.av_writeresponsevalid   ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                        //                .channel
		.rf_sink_ready           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_POSTED          (45),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.PKT_TRANS_LOCK            (48),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (50),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (79),
		.PKT_RESPONSE_STATUS_H     (87),
		.PKT_RESPONSE_STATUS_L     (86),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (88),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (89),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) apb_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (apb_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (apb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (apb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (apb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (apb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (apb_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (apb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (apb_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (apb_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (apb_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (apb_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (apb_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                             //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                             //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                              //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                       //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                           //                .channel
		.rf_sink_ready           (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (apb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (apb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50m_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50m_clk),                                                                           //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50m_clk),                                                                     //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (88),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                             //                .channel
		.rf_sink_ready           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) apb_m0_translator_avalon_universal_master_0_agent (
		.clk                     (syspll_c0_clk),                                                      //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.av_address              (apb_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (apb_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (apb_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (apb_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (apb_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (apb_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (apb_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (apb_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (apb_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (apb_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (apb_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (apb_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (apb_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (apb_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                          //          .ready
		.av_response             (),                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                                            //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                                            //                .valid
		.cp_data                 (crosser_002_out_data),                                                                             //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                                          //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_003_out_ready),                                                       //              cp.ready
		.cp_valid                (crosser_003_out_valid),                                                       //                .valid
		.cp_data                 (crosser_003_out_data),                                                        //                .data
		.cp_startofpacket        (crosser_003_out_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (crosser_003_out_endofpacket),                                                 //                .endofpacket
		.cp_channel              (crosser_003_out_channel),                                                     //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                 // (terminated)
		.csr_read          (1'b0),                                                                  // (terminated)
		.csr_write         (1'b0),                                                                  // (terminated)
		.csr_readdata      (),                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                  // (terminated)
		.almost_full_data  (),                                                                      // (terminated)
		.almost_empty_data (),                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                  // (terminated)
		.out_startofpacket (),                                                                      // (terminated)
		.out_endofpacket   (),                                                                      // (terminated)
		.in_empty          (1'b0),                                                                  // (terminated)
		.out_empty         (),                                                                      // (terminated)
		.in_error          (1'b0),                                                                  // (terminated)
		.out_error         (),                                                                      // (terminated)
		.in_channel        (1'b0),                                                                  // (terminated)
		.out_channel       ()                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_004_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_004_out_valid),                                                         //                .valid
		.cp_data                 (crosser_004_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_004_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_004_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_004_out_channel),                                                       //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_005_out_ready),                                                          //              cp.ready
		.cp_valid                (crosser_005_out_valid),                                                          //                .valid
		.cp_data                 (crosser_005_out_data),                                                           //                .data
		.cp_startofpacket        (crosser_005_out_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (crosser_005_out_endofpacket),                                                    //                .endofpacket
		.cp_channel              (crosser_005_out_channel),                                                        //                .channel
		.rf_sink_ready           (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.in_data           (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                    // (terminated)
		.csr_read          (1'b0),                                                                     // (terminated)
		.csr_write         (1'b0),                                                                     // (terminated)
		.csr_readdata      (),                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                     // (terminated)
		.almost_full_data  (),                                                                         // (terminated)
		.almost_empty_data (),                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                     // (terminated)
		.out_startofpacket (),                                                                         // (terminated)
		.out_endofpacket   (),                                                                         // (terminated)
		.in_empty          (1'b0),                                                                     // (terminated)
		.out_empty         (),                                                                         // (terminated)
		.in_error          (1'b0),                                                                     // (terminated)
		.out_error         (),                                                                         // (terminated)
		.in_channel        (1'b0),                                                                     // (terminated)
		.out_channel       ()                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                         //       clk_reset.reset
		.m0_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_006_out_ready),                                                      //              cp.ready
		.cp_valid                (crosser_006_out_valid),                                                      //                .valid
		.cp_data                 (crosser_006_out_data),                                                       //                .data
		.cp_startofpacket        (crosser_006_out_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (crosser_006_out_endofpacket),                                                //                .endofpacket
		.cp_channel              (crosser_006_out_channel),                                                    //                .channel
		.rf_sink_ready           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.in_data           (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                // (terminated)
		.csr_read          (1'b0),                                                                 // (terminated)
		.csr_write         (1'b0),                                                                 // (terminated)
		.csr_readdata      (),                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                 // (terminated)
		.almost_full_data  (),                                                                     // (terminated)
		.almost_empty_data (),                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                 // (terminated)
		.out_startofpacket (),                                                                     // (terminated)
		.out_endofpacket   (),                                                                     // (terminated)
		.in_empty          (1'b0),                                                                 // (terminated)
		.out_empty         (),                                                                     // (terminated)
		.in_error          (1'b0),                                                                 // (terminated)
		.out_error         (),                                                                     // (terminated)
		.in_channel        (1'b0),                                                                 // (terminated)
		.out_channel       ()                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_007_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_007_out_valid),                                                         //                .valid
		.cp_data                 (crosser_007_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_007_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_007_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_007_out_channel),                                                       //                .channel
		.rf_sink_ready           (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (hex_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) motora_duty_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (motora_duty_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_008_out_ready),                                                               //              cp.ready
		.cp_valid                (crosser_008_out_valid),                                                               //                .valid
		.cp_data                 (crosser_008_out_data),                                                                //                .data
		.cp_startofpacket        (crosser_008_out_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (crosser_008_out_endofpacket),                                                         //                .endofpacket
		.cp_channel              (crosser_008_out_channel),                                                             //                .channel
		.rf_sink_ready           (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (motora_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) motorb_duty_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (motorb_duty_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_009_out_ready),                                                               //              cp.ready
		.cp_valid                (crosser_009_out_valid),                                                               //                .valid
		.cp_data                 (crosser_009_out_data),                                                                //                .data
		.cp_startofpacket        (crosser_009_out_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (crosser_009_out_endofpacket),                                                         //                .endofpacket
		.cp_channel              (crosser_009_out_channel),                                                             //                .channel
		.rf_sink_ready           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) motora_dir_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (motora_dir_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_010_out_ready),                                                              //              cp.ready
		.cp_valid                (crosser_010_out_valid),                                                              //                .valid
		.cp_data                 (crosser_010_out_data),                                                               //                .data
		.cp_startofpacket        (crosser_010_out_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (crosser_010_out_endofpacket),                                                        //                .endofpacket
		.cp_channel              (crosser_010_out_channel),                                                            //                .channel
		.rf_sink_ready           (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (motora_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) motorb_dir_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (motorb_dir_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_011_out_ready),                                                              //              cp.ready
		.cp_valid                (crosser_011_out_valid),                                                              //                .valid
		.cp_data                 (crosser_011_out_data),                                                               //                .data
		.cp_startofpacket        (crosser_011_out_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (crosser_011_out_endofpacket),                                                        //                .endofpacket
		.cp_channel              (crosser_011_out_channel),                                                            //                .channel
		.rf_sink_ready           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_012_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_012_out_valid),                                                         //                .valid
		.cp_data                 (crosser_012_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_012_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_012_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_012_out_channel),                                                       //                .channel
		.rf_sink_ready           (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (hex_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) infra_sensor_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_013_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_013_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_013_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_013_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_013_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_013_out_channel),                                                                //                .channel
		.rf_sink_ready           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) infra_sensor_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_014_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_014_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_014_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_014_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_014_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_014_out_channel),                                                                //                .channel
		.rf_sink_ready           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) infra_sensor_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_015_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_015_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_015_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_015_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_015_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_015_out_channel),                                                                //                .channel
		.rf_sink_ready           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) infra_sensor_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_016_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_016_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_016_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_016_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_016_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_016_out_channel),                                                                //                .channel
		.rf_sink_ready           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) infra_sensor_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (syspll_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_017_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_017_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_017_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_017_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_017_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_017_out_channel),                                                                //                .channel
		.rf_sink_ready           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (syspll_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (syspll_c2_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	DE0Qsys_addr_router addr_router (
		.sink_ready         (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                                   //          .valid
		.src_data           (addr_router_src_data),                                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                              //          .endofpacket
	);

	DE0Qsys_addr_router_001 addr_router_001 (
		.sink_ready         (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                        //          .valid
		.src_data           (addr_router_001_src_data),                                                         //          .data
		.src_channel        (addr_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	DE0Qsys_addr_router_002 addr_router_002 (
		.sink_ready         (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                              //          .endofpacket
	);

	DE0Qsys_addr_router_002 addr_router_003 (
		.sink_ready         (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                    //          .valid
		.src_data           (addr_router_003_src_data),                                                     //          .data
		.src_channel        (addr_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                               //          .endofpacket
	);

	DE0Qsys_id_router id_router (
		.sink_ready         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	DE0Qsys_id_router_001 id_router_001 (
		.sink_ready         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_ctrl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	DE0Qsys_id_router_002 id_router_002 (
		.sink_ready         (apb_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (apb_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (apb_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (apb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (apb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                           //          .valid
		.src_data           (id_router_002_src_data),                                            //          .data
		.src_channel        (id_router_002_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                      //          .endofpacket
	);

	DE0Qsys_id_router_003 id_router_003 (
		.sink_ready         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (syspll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50m_clk),                                                                 //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                     //       src.ready
		.src_valid          (id_router_003_src_valid),                                                     //          .valid
		.src_data           (id_router_003_src_data),                                                      //          .data
		.src_channel        (id_router_003_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                //          .endofpacket
	);

	DE0Qsys_id_router_003 id_router_004 (
		.sink_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                           //       src.ready
		.src_valid          (id_router_004_src_valid),                                                           //          .valid
		.src_data           (id_router_004_src_data),                                                            //          .data
		.src_channel        (id_router_004_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                      //          .endofpacket
	);

	DE0Qsys_addr_router_004 addr_router_004 (
		.sink_ready         (apb_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (apb_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (apb_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (apb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (apb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (syspll_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                          //       src.ready
		.src_valid          (addr_router_004_src_valid),                                          //          .valid
		.src_data           (addr_router_004_src_data),                                           //          .data
		.src_channel        (addr_router_004_src_channel),                                        //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                     //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_006 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                           //       src.ready
		.src_valid          (id_router_006_src_valid),                                           //          .valid
		.src_data           (id_router_006_src_data),                                            //          .data
		.src_channel        (id_router_006_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                      //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_007 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                             //       src.ready
		.src_valid          (id_router_007_src_valid),                                             //          .valid
		.src_data           (id_router_007_src_data),                                              //          .data
		.src_channel        (id_router_007_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                        //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_008 (
		.sink_ready         (button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                              //       src.ready
		.src_valid          (id_router_008_src_valid),                                              //          .valid
		.src_data           (id_router_008_src_data),                                               //          .data
		.src_channel        (id_router_008_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                         //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_009 (
		.sink_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                               // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                          //       src.ready
		.src_valid          (id_router_009_src_valid),                                          //          .valid
		.src_data           (id_router_009_src_data),                                           //          .data
		.src_channel        (id_router_009_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                     //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_010 (
		.sink_ready         (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                             //       src.ready
		.src_valid          (id_router_010_src_valid),                                             //          .valid
		.src_data           (id_router_010_src_data),                                              //          .data
		.src_channel        (id_router_010_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                        //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_011 (
		.sink_ready         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (motora_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                   //       src.ready
		.src_valid          (id_router_011_src_valid),                                                   //          .valid
		.src_data           (id_router_011_src_data),                                                    //          .data
		.src_channel        (id_router_011_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                              //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_012 (
		.sink_ready         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (motorb_duty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                   //       src.ready
		.src_valid          (id_router_012_src_valid),                                                   //          .valid
		.src_data           (id_router_012_src_data),                                                    //          .data
		.src_channel        (id_router_012_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                              //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_013 (
		.sink_ready         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (motora_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_014 (
		.sink_ready         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (motorb_dir_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                             //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_015 (
		.sink_ready         (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                             //       src.ready
		.src_valid          (id_router_015_src_valid),                                             //          .valid
		.src_data           (id_router_015_src_data),                                              //          .data
		.src_channel        (id_router_015_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                        //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_016 (
		.sink_ready         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (infra_sensor_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                      //       src.ready
		.src_valid          (id_router_016_src_valid),                                                      //          .valid
		.src_data           (id_router_016_src_data),                                                       //          .data
		.src_channel        (id_router_016_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                 //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_017 (
		.sink_ready         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (infra_sensor_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                      //       src.ready
		.src_valid          (id_router_017_src_valid),                                                      //          .valid
		.src_data           (id_router_017_src_data),                                                       //          .data
		.src_channel        (id_router_017_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                 //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_018 (
		.sink_ready         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (infra_sensor_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                      //       src.ready
		.src_valid          (id_router_018_src_valid),                                                      //          .valid
		.src_data           (id_router_018_src_data),                                                       //          .data
		.src_channel        (id_router_018_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                 //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_019 (
		.sink_ready         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (infra_sensor_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                      //       src.ready
		.src_valid          (id_router_019_src_valid),                                                      //          .valid
		.src_data           (id_router_019_src_data),                                                       //          .data
		.src_channel        (id_router_019_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                 //          .endofpacket
	);

	DE0Qsys_id_router_005 id_router_020 (
		.sink_ready         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (infra_sensor_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (syspll_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                      //       src.ready
		.src_valid          (id_router_020_src_valid),                                                      //          .valid
		.src_data           (id_router_020_src_data),                                                       //          .data
		.src_channel        (id_router_020_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                 //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.VALID_WIDTH               (5),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (syspll_c0_clk),                      //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (16),
		.VALID_WIDTH               (16),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (syspll_c0_clk),                      //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_004_src_data),           //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_004_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_004_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_004_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (70),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (50),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.PKT_BURST_TYPE_H          (67),
		.PKT_BURST_TYPE_L          (66),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (88),
		.ST_CHANNEL_W              (5),
		.OUT_BYTE_CNT_H            (51),
		.OUT_BURSTWRAP_H           (62),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (syspll_c0_clk),                       //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (88),
		.PKT_BYTE_CNT_H            (77),
		.PKT_BYTE_CNT_L            (68),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (78),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (5),
		.OUT_BYTE_CNT_H            (70),
		.OUT_BURSTWRAP_H           (80),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (syspll_c0_clk),                           //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (nios2cpu_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                         // reset_in1.reset
		.clk        (syspll_c0_clk),                          //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                       // (terminated)
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                         // reset_in0.reset
		.reset_in1  (nios2cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (syspll_c2_clk),                          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req  (),                                       // (terminated)
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_50m_clk),                        //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	DE0Qsys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (syspll_c0_clk),                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (syspll_c0_clk),                         //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                 //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),               //           .channel
		.sink_data          (limiter_cmd_src_data),                  //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),         //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),           //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)    //           .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_mux_001 cmd_xbar_mux_002 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_003 rsp_xbar_demux (
		.clk                (syspll_c0_clk),                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_001 rsp_xbar_demux_002 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_50m_clk),                           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (syspll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (crosser_001_out_ready),                 //     sink3.ready
		.sink3_valid         (crosser_001_out_valid),                 //          .valid
		.sink3_channel       (crosser_001_out_channel),               //          .channel
		.sink3_data          (crosser_001_out_data),                  //          .data
		.sink3_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink3_endofpacket   (crosser_001_out_endofpacket),           //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_002_src2_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_002_src2_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_002 rsp_xbar_mux_003 (
		.clk                 (syspll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_002_src3_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	DE0Qsys_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                 (syspll_c0_clk),                          //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_004_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_004_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_004_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_004_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_004_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_004_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_004_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_004_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_004_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_004_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_004_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_004_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_004_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_004_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_004_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_004_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_004_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_004_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_004_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_004_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_004_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_004_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_004_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_004_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_004_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_004_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_004_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_004_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_004_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_004_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_004_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_004_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_004_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_004_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_004_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_004_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_004_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_004_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_004_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_004_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_004_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_004_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_004_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_004_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_004_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_004_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_004_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_004_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_004_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_004_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_004_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_004_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_004_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_004_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_004_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_004_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_004_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_004_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_004_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_004_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_004_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_004_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_004_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_004_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_004_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_004_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_004_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_004_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_004_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_004_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_004_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_004_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_004_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_004_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_004_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_004_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_004_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_004_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_004_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_004_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_004_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_004_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_004_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_004_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_004_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_004_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_004_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_004_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_004_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_004_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_004_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_004_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_004_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_004_src15_endofpacket)    //           .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_007 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_008 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_009 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_012 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_013 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_014 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_015 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_016 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_017 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_018 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_019 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_demux_005 rsp_xbar_demux_020 (
		.clk                (syspll_c2_clk),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	DE0Qsys_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                  (syspll_c0_clk),                      //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.src_ready            (rsp_xbar_mux_004_src_ready),         //       src.ready
		.src_valid            (rsp_xbar_mux_004_src_valid),         //          .valid
		.src_data             (rsp_xbar_mux_004_src_data),          //          .data
		.src_channel          (rsp_xbar_mux_004_src_channel),       //          .channel
		.src_startofpacket    (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.sink0_ready          (crosser_018_out_ready),              //     sink0.ready
		.sink0_valid          (crosser_018_out_valid),              //          .valid
		.sink0_channel        (crosser_018_out_channel),            //          .channel
		.sink0_data           (crosser_018_out_data),               //          .data
		.sink0_startofpacket  (crosser_018_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket    (crosser_018_out_endofpacket),        //          .endofpacket
		.sink1_ready          (crosser_019_out_ready),              //     sink1.ready
		.sink1_valid          (crosser_019_out_valid),              //          .valid
		.sink1_channel        (crosser_019_out_channel),            //          .channel
		.sink1_data           (crosser_019_out_data),               //          .data
		.sink1_startofpacket  (crosser_019_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket    (crosser_019_out_endofpacket),        //          .endofpacket
		.sink2_ready          (crosser_020_out_ready),              //     sink2.ready
		.sink2_valid          (crosser_020_out_valid),              //          .valid
		.sink2_channel        (crosser_020_out_channel),            //          .channel
		.sink2_data           (crosser_020_out_data),               //          .data
		.sink2_startofpacket  (crosser_020_out_startofpacket),      //          .startofpacket
		.sink2_endofpacket    (crosser_020_out_endofpacket),        //          .endofpacket
		.sink3_ready          (crosser_021_out_ready),              //     sink3.ready
		.sink3_valid          (crosser_021_out_valid),              //          .valid
		.sink3_channel        (crosser_021_out_channel),            //          .channel
		.sink3_data           (crosser_021_out_data),               //          .data
		.sink3_startofpacket  (crosser_021_out_startofpacket),      //          .startofpacket
		.sink3_endofpacket    (crosser_021_out_endofpacket),        //          .endofpacket
		.sink4_ready          (crosser_022_out_ready),              //     sink4.ready
		.sink4_valid          (crosser_022_out_valid),              //          .valid
		.sink4_channel        (crosser_022_out_channel),            //          .channel
		.sink4_data           (crosser_022_out_data),               //          .data
		.sink4_startofpacket  (crosser_022_out_startofpacket),      //          .startofpacket
		.sink4_endofpacket    (crosser_022_out_endofpacket),        //          .endofpacket
		.sink5_ready          (crosser_023_out_ready),              //     sink5.ready
		.sink5_valid          (crosser_023_out_valid),              //          .valid
		.sink5_channel        (crosser_023_out_channel),            //          .channel
		.sink5_data           (crosser_023_out_data),               //          .data
		.sink5_startofpacket  (crosser_023_out_startofpacket),      //          .startofpacket
		.sink5_endofpacket    (crosser_023_out_endofpacket),        //          .endofpacket
		.sink6_ready          (crosser_024_out_ready),              //     sink6.ready
		.sink6_valid          (crosser_024_out_valid),              //          .valid
		.sink6_channel        (crosser_024_out_channel),            //          .channel
		.sink6_data           (crosser_024_out_data),               //          .data
		.sink6_startofpacket  (crosser_024_out_startofpacket),      //          .startofpacket
		.sink6_endofpacket    (crosser_024_out_endofpacket),        //          .endofpacket
		.sink7_ready          (crosser_025_out_ready),              //     sink7.ready
		.sink7_valid          (crosser_025_out_valid),              //          .valid
		.sink7_channel        (crosser_025_out_channel),            //          .channel
		.sink7_data           (crosser_025_out_data),               //          .data
		.sink7_startofpacket  (crosser_025_out_startofpacket),      //          .startofpacket
		.sink7_endofpacket    (crosser_025_out_endofpacket),        //          .endofpacket
		.sink8_ready          (crosser_026_out_ready),              //     sink8.ready
		.sink8_valid          (crosser_026_out_valid),              //          .valid
		.sink8_channel        (crosser_026_out_channel),            //          .channel
		.sink8_data           (crosser_026_out_data),               //          .data
		.sink8_startofpacket  (crosser_026_out_startofpacket),      //          .startofpacket
		.sink8_endofpacket    (crosser_026_out_endofpacket),        //          .endofpacket
		.sink9_ready          (crosser_027_out_ready),              //     sink9.ready
		.sink9_valid          (crosser_027_out_valid),              //          .valid
		.sink9_channel        (crosser_027_out_channel),            //          .channel
		.sink9_data           (crosser_027_out_data),               //          .data
		.sink9_startofpacket  (crosser_027_out_startofpacket),      //          .startofpacket
		.sink9_endofpacket    (crosser_027_out_endofpacket),        //          .endofpacket
		.sink10_ready         (crosser_028_out_ready),              //    sink10.ready
		.sink10_valid         (crosser_028_out_valid),              //          .valid
		.sink10_channel       (crosser_028_out_channel),            //          .channel
		.sink10_data          (crosser_028_out_data),               //          .data
		.sink10_startofpacket (crosser_028_out_startofpacket),      //          .startofpacket
		.sink10_endofpacket   (crosser_028_out_endofpacket),        //          .endofpacket
		.sink11_ready         (crosser_029_out_ready),              //    sink11.ready
		.sink11_valid         (crosser_029_out_valid),              //          .valid
		.sink11_channel       (crosser_029_out_channel),            //          .channel
		.sink11_data          (crosser_029_out_data),               //          .data
		.sink11_startofpacket (crosser_029_out_startofpacket),      //          .startofpacket
		.sink11_endofpacket   (crosser_029_out_endofpacket),        //          .endofpacket
		.sink12_ready         (crosser_030_out_ready),              //    sink12.ready
		.sink12_valid         (crosser_030_out_valid),              //          .valid
		.sink12_channel       (crosser_030_out_channel),            //          .channel
		.sink12_data          (crosser_030_out_data),               //          .data
		.sink12_startofpacket (crosser_030_out_startofpacket),      //          .startofpacket
		.sink12_endofpacket   (crosser_030_out_endofpacket),        //          .endofpacket
		.sink13_ready         (crosser_031_out_ready),              //    sink13.ready
		.sink13_valid         (crosser_031_out_valid),              //          .valid
		.sink13_channel       (crosser_031_out_channel),            //          .channel
		.sink13_data          (crosser_031_out_data),               //          .data
		.sink13_startofpacket (crosser_031_out_startofpacket),      //          .startofpacket
		.sink13_endofpacket   (crosser_031_out_endofpacket),        //          .endofpacket
		.sink14_ready         (crosser_032_out_ready),              //    sink14.ready
		.sink14_valid         (crosser_032_out_valid),              //          .valid
		.sink14_channel       (crosser_032_out_channel),            //          .channel
		.sink14_data          (crosser_032_out_data),               //          .data
		.sink14_startofpacket (crosser_032_out_startofpacket),      //          .startofpacket
		.sink14_endofpacket   (crosser_032_out_endofpacket),        //          .endofpacket
		.sink15_ready         (crosser_033_out_ready),              //    sink15.ready
		.sink15_valid         (crosser_033_out_valid),              //          .valid
		.sink15_channel       (crosser_033_out_channel),            //          .channel
		.sink15_data          (crosser_033_out_data),               //          .data
		.sink15_startofpacket (crosser_033_out_startofpacket),      //          .startofpacket
		.sink15_endofpacket   (crosser_033_out_endofpacket)         //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (61),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (77),
		.IN_PKT_BYTE_CNT_L             (68),
		.IN_PKT_TRANS_COMPRESSED_READ  (62),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (78),
		.IN_PKT_BURST_SIZE_H           (83),
		.IN_PKT_BURST_SIZE_L           (81),
		.IN_PKT_RESPONSE_STATUS_H      (105),
		.IN_PKT_RESPONSE_STATUS_L      (104),
		.IN_PKT_TRANS_EXCLUSIVE        (67),
		.IN_PKT_BURST_TYPE_H           (85),
		.IN_PKT_BURST_TYPE_L           (84),
		.IN_ST_DATA_W                  (106),
		.OUT_PKT_ADDR_H                (43),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (59),
		.OUT_PKT_BYTE_CNT_L            (50),
		.OUT_PKT_TRANS_COMPRESSED_READ (44),
		.OUT_PKT_BURST_SIZE_H          (65),
		.OUT_PKT_BURST_SIZE_L          (63),
		.OUT_PKT_RESPONSE_STATUS_H     (87),
		.OUT_PKT_RESPONSE_STATUS_L     (86),
		.OUT_PKT_TRANS_EXCLUSIVE       (49),
		.OUT_PKT_BURST_TYPE_H          (67),
		.OUT_PKT_BURST_TYPE_L          (66),
		.OUT_ST_DATA_W                 (88),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (syspll_c0_clk),                      //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (43),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (59),
		.IN_PKT_BYTE_CNT_L             (50),
		.IN_PKT_TRANS_COMPRESSED_READ  (44),
		.IN_PKT_BURSTWRAP_H            (62),
		.IN_PKT_BURSTWRAP_L            (60),
		.IN_PKT_BURST_SIZE_H           (65),
		.IN_PKT_BURST_SIZE_L           (63),
		.IN_PKT_RESPONSE_STATUS_H      (87),
		.IN_PKT_RESPONSE_STATUS_L      (86),
		.IN_PKT_TRANS_EXCLUSIVE        (49),
		.IN_PKT_BURST_TYPE_H           (67),
		.IN_PKT_BURST_TYPE_L           (66),
		.IN_ST_DATA_W                  (88),
		.OUT_PKT_ADDR_H                (61),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (77),
		.OUT_PKT_BYTE_CNT_L            (68),
		.OUT_PKT_TRANS_COMPRESSED_READ (62),
		.OUT_PKT_BURST_SIZE_H          (83),
		.OUT_PKT_BURST_SIZE_L          (81),
		.OUT_PKT_RESPONSE_STATUS_H     (105),
		.OUT_PKT_RESPONSE_STATUS_L     (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (67),
		.OUT_PKT_BURST_TYPE_H          (85),
		.OUT_PKT_BURST_TYPE_L          (84),
		.OUT_ST_DATA_W                 (106),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (syspll_c0_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (106),
		.BITS_PER_SYMBOL     (106),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (5),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_50m_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src3_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src3_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src3_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src3_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src3_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (106),
		.BITS_PER_SYMBOL     (106),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (5),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_50m_clk),                           //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_003_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_003_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_003_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_003_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src1_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src1_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src1_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src1_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src2_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src2_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src2_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src2_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src2_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src2_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src3_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src3_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src3_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src3_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src3_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src3_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src4_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src5_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src6_data),          //              .data
		.out_ready         (crosser_008_out_ready),                 //           out.ready
		.out_valid         (crosser_008_out_valid),                 //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_008_out_channel),               //              .channel
		.out_data          (crosser_008_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src7_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src7_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src7_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src7_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src7_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src7_data),          //              .data
		.out_ready         (crosser_009_out_ready),                 //           out.ready
		.out_valid         (crosser_009_out_valid),                 //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_009_out_channel),               //              .channel
		.out_data          (crosser_009_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_010 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src8_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src8_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src8_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src8_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src8_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src8_data),          //              .data
		.out_ready         (crosser_010_out_ready),                 //           out.ready
		.out_valid         (crosser_010_out_valid),                 //              .valid
		.out_startofpacket (crosser_010_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_010_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_010_out_channel),               //              .channel
		.out_data          (crosser_010_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_011 (
		.in_clk            (syspll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src9_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src9_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src9_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src9_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src9_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src9_data),          //              .data
		.out_ready         (crosser_011_out_ready),                 //           out.ready
		.out_valid         (crosser_011_out_valid),                 //              .valid
		.out_startofpacket (crosser_011_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_011_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_011_out_channel),               //              .channel
		.out_data          (crosser_011_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_012 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src10_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src10_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src10_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src10_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src10_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src10_data),          //              .data
		.out_ready         (crosser_012_out_ready),                  //           out.ready
		.out_valid         (crosser_012_out_valid),                  //              .valid
		.out_startofpacket (crosser_012_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_012_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_012_out_channel),                //              .channel
		.out_data          (crosser_012_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_013 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src11_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src11_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src11_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src11_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src11_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src11_data),          //              .data
		.out_ready         (crosser_013_out_ready),                  //           out.ready
		.out_valid         (crosser_013_out_valid),                  //              .valid
		.out_startofpacket (crosser_013_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_013_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_013_out_channel),                //              .channel
		.out_data          (crosser_013_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_014 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src12_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src12_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src12_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src12_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src12_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src12_data),          //              .data
		.out_ready         (crosser_014_out_ready),                  //           out.ready
		.out_valid         (crosser_014_out_valid),                  //              .valid
		.out_startofpacket (crosser_014_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_014_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_014_out_channel),                //              .channel
		.out_data          (crosser_014_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_015 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src13_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src13_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src13_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src13_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src13_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src13_data),          //              .data
		.out_ready         (crosser_015_out_ready),                  //           out.ready
		.out_valid         (crosser_015_out_valid),                  //              .valid
		.out_startofpacket (crosser_015_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_015_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_015_out_channel),                //              .channel
		.out_data          (crosser_015_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_016 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src14_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src14_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src14_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src14_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src14_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src14_data),          //              .data
		.out_ready         (crosser_016_out_ready),                  //           out.ready
		.out_valid         (crosser_016_out_valid),                  //              .valid
		.out_startofpacket (crosser_016_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_016_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_016_out_channel),                //              .channel
		.out_data          (crosser_016_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_017 (
		.in_clk            (syspll_c0_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (syspll_c2_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src15_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src15_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src15_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src15_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src15_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src15_data),          //              .data
		.out_ready         (crosser_017_out_ready),                  //           out.ready
		.out_valid         (crosser_017_out_valid),                  //              .valid
		.out_startofpacket (crosser_017_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_017_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_017_out_channel),                //              .channel
		.out_data          (crosser_017_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_018 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_018_out_ready),                 //           out.ready
		.out_valid         (crosser_018_out_valid),                 //              .valid
		.out_startofpacket (crosser_018_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_018_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_018_out_channel),               //              .channel
		.out_data          (crosser_018_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_019 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_019_out_ready),                 //           out.ready
		.out_valid         (crosser_019_out_valid),                 //              .valid
		.out_startofpacket (crosser_019_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_019_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_019_out_channel),               //              .channel
		.out_data          (crosser_019_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_020 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_020_out_ready),                 //           out.ready
		.out_valid         (crosser_020_out_valid),                 //              .valid
		.out_startofpacket (crosser_020_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_020_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_020_out_channel),               //              .channel
		.out_data          (crosser_020_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_021 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_021_out_ready),                 //           out.ready
		.out_valid         (crosser_021_out_valid),                 //              .valid
		.out_startofpacket (crosser_021_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_021_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_021_out_channel),               //              .channel
		.out_data          (crosser_021_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_022 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_009_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_009_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_009_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_009_src0_data),          //              .data
		.out_ready         (crosser_022_out_ready),                 //           out.ready
		.out_valid         (crosser_022_out_valid),                 //              .valid
		.out_startofpacket (crosser_022_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_022_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_022_out_channel),               //              .channel
		.out_data          (crosser_022_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_023 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_010_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_010_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_010_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_010_src0_data),          //              .data
		.out_ready         (crosser_023_out_ready),                 //           out.ready
		.out_valid         (crosser_023_out_valid),                 //              .valid
		.out_startofpacket (crosser_023_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_023_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_023_out_channel),               //              .channel
		.out_data          (crosser_023_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_024 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_011_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_011_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_011_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_011_src0_data),          //              .data
		.out_ready         (crosser_024_out_ready),                 //           out.ready
		.out_valid         (crosser_024_out_valid),                 //              .valid
		.out_startofpacket (crosser_024_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_024_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_024_out_channel),               //              .channel
		.out_data          (crosser_024_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_025 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_025_out_ready),                 //           out.ready
		.out_valid         (crosser_025_out_valid),                 //              .valid
		.out_startofpacket (crosser_025_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_025_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_025_out_channel),               //              .channel
		.out_data          (crosser_025_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_026 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_026_out_ready),                 //           out.ready
		.out_valid         (crosser_026_out_valid),                 //              .valid
		.out_startofpacket (crosser_026_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_026_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_026_out_channel),               //              .channel
		.out_data          (crosser_026_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_027 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_014_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_014_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_014_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_014_src0_data),          //              .data
		.out_ready         (crosser_027_out_ready),                 //           out.ready
		.out_valid         (crosser_027_out_valid),                 //              .valid
		.out_startofpacket (crosser_027_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_027_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_027_out_channel),               //              .channel
		.out_data          (crosser_027_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_028 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_015_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_015_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_015_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_015_src0_data),          //              .data
		.out_ready         (crosser_028_out_ready),                 //           out.ready
		.out_valid         (crosser_028_out_valid),                 //              .valid
		.out_startofpacket (crosser_028_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_028_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_028_out_channel),               //              .channel
		.out_data          (crosser_028_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_029 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_016_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_016_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_016_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_016_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_016_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_016_src0_data),          //              .data
		.out_ready         (crosser_029_out_ready),                 //           out.ready
		.out_valid         (crosser_029_out_valid),                 //              .valid
		.out_startofpacket (crosser_029_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_029_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_029_out_channel),               //              .channel
		.out_data          (crosser_029_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_030 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_017_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_017_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_017_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_017_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_017_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_017_src0_data),          //              .data
		.out_ready         (crosser_030_out_ready),                 //           out.ready
		.out_valid         (crosser_030_out_valid),                 //              .valid
		.out_startofpacket (crosser_030_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_030_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_030_out_channel),               //              .channel
		.out_data          (crosser_030_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_031 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_018_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_018_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_018_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_018_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_018_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_018_src0_data),          //              .data
		.out_ready         (crosser_031_out_ready),                 //           out.ready
		.out_valid         (crosser_031_out_valid),                 //              .valid
		.out_startofpacket (crosser_031_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_031_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_031_out_channel),               //              .channel
		.out_data          (crosser_031_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_032 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_019_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_019_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_019_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_019_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_019_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_019_src0_data),          //              .data
		.out_ready         (crosser_032_out_ready),                 //           out.ready
		.out_valid         (crosser_032_out_valid),                 //              .valid
		.out_startofpacket (crosser_032_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_032_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_032_out_channel),               //              .channel
		.out_data          (crosser_032_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_033 (
		.in_clk            (syspll_c2_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (syspll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_020_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_020_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_020_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_020_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_020_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_020_src0_data),          //              .data
		.out_ready         (crosser_033_out_ready),                 //           out.ready
		.out_valid         (crosser_033_out_valid),                 //              .valid
		.out_startofpacket (crosser_033_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_033_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_033_out_channel),               //              .channel
		.out_data          (crosser_033_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	DE0Qsys_irq_mapper irq_mapper (
		.clk           (syspll_c0_clk),                  //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2cpu_d_irq_irq)              //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (syspll_c2_clk),                      //       receiver_clk.clk
		.sender_clk     (syspll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (syspll_c2_clk),                      //       receiver_clk.clk
		.sender_clk     (syspll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

endmodule
